magic
tech sky130A
magscale 1 2
timestamp 1712109191
<< nwell >>
rect -2290 -797 2290 797
<< mvpmos >>
rect -2032 -500 -1632 500
rect -1574 -500 -1174 500
rect -1116 -500 -716 500
rect -658 -500 -258 500
rect -200 -500 200 500
rect 258 -500 658 500
rect 716 -500 1116 500
rect 1174 -500 1574 500
rect 1632 -500 2032 500
<< mvpdiff >>
rect -2090 488 -2032 500
rect -2090 -488 -2078 488
rect -2044 -488 -2032 488
rect -2090 -500 -2032 -488
rect -1632 488 -1574 500
rect -1632 -488 -1620 488
rect -1586 -488 -1574 488
rect -1632 -500 -1574 -488
rect -1174 488 -1116 500
rect -1174 -488 -1162 488
rect -1128 -488 -1116 488
rect -1174 -500 -1116 -488
rect -716 488 -658 500
rect -716 -488 -704 488
rect -670 -488 -658 488
rect -716 -500 -658 -488
rect -258 488 -200 500
rect -258 -488 -246 488
rect -212 -488 -200 488
rect -258 -500 -200 -488
rect 200 488 258 500
rect 200 -488 212 488
rect 246 -488 258 488
rect 200 -500 258 -488
rect 658 488 716 500
rect 658 -488 670 488
rect 704 -488 716 488
rect 658 -500 716 -488
rect 1116 488 1174 500
rect 1116 -488 1128 488
rect 1162 -488 1174 488
rect 1116 -500 1174 -488
rect 1574 488 1632 500
rect 1574 -488 1586 488
rect 1620 -488 1632 488
rect 1574 -500 1632 -488
rect 2032 488 2090 500
rect 2032 -488 2044 488
rect 2078 -488 2090 488
rect 2032 -500 2090 -488
<< mvpdiffc >>
rect -2078 -488 -2044 488
rect -1620 -488 -1586 488
rect -1162 -488 -1128 488
rect -704 -488 -670 488
rect -246 -488 -212 488
rect 212 -488 246 488
rect 670 -488 704 488
rect 1128 -488 1162 488
rect 1586 -488 1620 488
rect 2044 -488 2078 488
<< mvnsubdiff >>
rect -2224 719 2224 731
rect -2224 685 -2116 719
rect 2116 685 2224 719
rect -2224 673 2224 685
rect -2224 623 -2166 673
rect -2224 -623 -2212 623
rect -2178 -623 -2166 623
rect 2166 623 2224 673
rect -2224 -673 -2166 -623
rect 2166 -623 2178 623
rect 2212 -623 2224 623
rect 2166 -673 2224 -623
rect -2224 -685 2224 -673
rect -2224 -719 -2116 -685
rect 2116 -719 2224 -685
rect -2224 -731 2224 -719
<< mvnsubdiffcont >>
rect -2116 685 2116 719
rect -2212 -623 -2178 623
rect 2178 -623 2212 623
rect -2116 -719 2116 -685
<< poly >>
rect -2032 581 -1632 597
rect -2032 547 -2016 581
rect -1648 547 -1632 581
rect -2032 500 -1632 547
rect -1574 581 -1174 597
rect -1574 547 -1558 581
rect -1190 547 -1174 581
rect -1574 500 -1174 547
rect -1116 581 -716 597
rect -1116 547 -1100 581
rect -732 547 -716 581
rect -1116 500 -716 547
rect -658 581 -258 597
rect -658 547 -642 581
rect -274 547 -258 581
rect -658 500 -258 547
rect -200 581 200 597
rect -200 547 -184 581
rect 184 547 200 581
rect -200 500 200 547
rect 258 581 658 597
rect 258 547 274 581
rect 642 547 658 581
rect 258 500 658 547
rect 716 581 1116 597
rect 716 547 732 581
rect 1100 547 1116 581
rect 716 500 1116 547
rect 1174 581 1574 597
rect 1174 547 1190 581
rect 1558 547 1574 581
rect 1174 500 1574 547
rect 1632 581 2032 597
rect 1632 547 1648 581
rect 2016 547 2032 581
rect 1632 500 2032 547
rect -2032 -547 -1632 -500
rect -2032 -581 -2016 -547
rect -1648 -581 -1632 -547
rect -2032 -597 -1632 -581
rect -1574 -547 -1174 -500
rect -1574 -581 -1558 -547
rect -1190 -581 -1174 -547
rect -1574 -597 -1174 -581
rect -1116 -547 -716 -500
rect -1116 -581 -1100 -547
rect -732 -581 -716 -547
rect -1116 -597 -716 -581
rect -658 -547 -258 -500
rect -658 -581 -642 -547
rect -274 -581 -258 -547
rect -658 -597 -258 -581
rect -200 -547 200 -500
rect -200 -581 -184 -547
rect 184 -581 200 -547
rect -200 -597 200 -581
rect 258 -547 658 -500
rect 258 -581 274 -547
rect 642 -581 658 -547
rect 258 -597 658 -581
rect 716 -547 1116 -500
rect 716 -581 732 -547
rect 1100 -581 1116 -547
rect 716 -597 1116 -581
rect 1174 -547 1574 -500
rect 1174 -581 1190 -547
rect 1558 -581 1574 -547
rect 1174 -597 1574 -581
rect 1632 -547 2032 -500
rect 1632 -581 1648 -547
rect 2016 -581 2032 -547
rect 1632 -597 2032 -581
<< polycont >>
rect -2016 547 -1648 581
rect -1558 547 -1190 581
rect -1100 547 -732 581
rect -642 547 -274 581
rect -184 547 184 581
rect 274 547 642 581
rect 732 547 1100 581
rect 1190 547 1558 581
rect 1648 547 2016 581
rect -2016 -581 -1648 -547
rect -1558 -581 -1190 -547
rect -1100 -581 -732 -547
rect -642 -581 -274 -547
rect -184 -581 184 -547
rect 274 -581 642 -547
rect 732 -581 1100 -547
rect 1190 -581 1558 -547
rect 1648 -581 2016 -547
<< locali >>
rect -2212 685 -2116 719
rect 2116 685 2212 719
rect -2212 623 -2178 685
rect 2178 623 2212 685
rect -2032 547 -2016 581
rect -1648 547 -1632 581
rect -1574 547 -1558 581
rect -1190 547 -1174 581
rect -1116 547 -1100 581
rect -732 547 -716 581
rect -658 547 -642 581
rect -274 547 -258 581
rect -200 547 -184 581
rect 184 547 200 581
rect 258 547 274 581
rect 642 547 658 581
rect 716 547 732 581
rect 1100 547 1116 581
rect 1174 547 1190 581
rect 1558 547 1574 581
rect 1632 547 1648 581
rect 2016 547 2032 581
rect -2078 488 -2044 504
rect -2078 -504 -2044 -488
rect -1620 488 -1586 504
rect -1620 -504 -1586 -488
rect -1162 488 -1128 504
rect -1162 -504 -1128 -488
rect -704 488 -670 504
rect -704 -504 -670 -488
rect -246 488 -212 504
rect -246 -504 -212 -488
rect 212 488 246 504
rect 212 -504 246 -488
rect 670 488 704 504
rect 670 -504 704 -488
rect 1128 488 1162 504
rect 1128 -504 1162 -488
rect 1586 488 1620 504
rect 1586 -504 1620 -488
rect 2044 488 2078 504
rect 2044 -504 2078 -488
rect -2032 -581 -2016 -547
rect -1648 -581 -1632 -547
rect -1574 -581 -1558 -547
rect -1190 -581 -1174 -547
rect -1116 -581 -1100 -547
rect -732 -581 -716 -547
rect -658 -581 -642 -547
rect -274 -581 -258 -547
rect -200 -581 -184 -547
rect 184 -581 200 -547
rect 258 -581 274 -547
rect 642 -581 658 -547
rect 716 -581 732 -547
rect 1100 -581 1116 -547
rect 1174 -581 1190 -547
rect 1558 -581 1574 -547
rect 1632 -581 1648 -547
rect 2016 -581 2032 -547
rect -2212 -685 -2178 -623
rect 2178 -685 2212 -623
rect -2212 -719 -2116 -685
rect 2116 -719 2212 -685
<< viali >>
rect -2016 547 -1648 581
rect -1558 547 -1190 581
rect -1100 547 -732 581
rect -642 547 -274 581
rect -184 547 184 581
rect 274 547 642 581
rect 732 547 1100 581
rect 1190 547 1558 581
rect 1648 547 2016 581
rect -2078 -488 -2044 488
rect -1620 -488 -1586 488
rect -1162 -488 -1128 488
rect -704 -488 -670 488
rect -246 -488 -212 488
rect 212 -488 246 488
rect 670 -488 704 488
rect 1128 -488 1162 488
rect 1586 -488 1620 488
rect 2044 -488 2078 488
rect -2016 -581 -1648 -547
rect -1558 -581 -1190 -547
rect -1100 -581 -732 -547
rect -642 -581 -274 -547
rect -184 -581 184 -547
rect 274 -581 642 -547
rect 732 -581 1100 -547
rect 1190 -581 1558 -547
rect 1648 -581 2016 -547
<< metal1 >>
rect -2028 581 -1636 587
rect -2028 547 -2016 581
rect -1648 547 -1636 581
rect -2028 541 -1636 547
rect -1570 581 -1178 587
rect -1570 547 -1558 581
rect -1190 547 -1178 581
rect -1570 541 -1178 547
rect -1112 581 -720 587
rect -1112 547 -1100 581
rect -732 547 -720 581
rect -1112 541 -720 547
rect -654 581 -262 587
rect -654 547 -642 581
rect -274 547 -262 581
rect -654 541 -262 547
rect -196 581 196 587
rect -196 547 -184 581
rect 184 547 196 581
rect -196 541 196 547
rect 262 581 654 587
rect 262 547 274 581
rect 642 547 654 581
rect 262 541 654 547
rect 720 581 1112 587
rect 720 547 732 581
rect 1100 547 1112 581
rect 720 541 1112 547
rect 1178 581 1570 587
rect 1178 547 1190 581
rect 1558 547 1570 581
rect 1178 541 1570 547
rect 1636 581 2028 587
rect 1636 547 1648 581
rect 2016 547 2028 581
rect 1636 541 2028 547
rect -2084 488 -2038 500
rect -2084 -488 -2078 488
rect -2044 -488 -2038 488
rect -2084 -500 -2038 -488
rect -1626 488 -1580 500
rect -1626 -488 -1620 488
rect -1586 -488 -1580 488
rect -1626 -500 -1580 -488
rect -1168 488 -1122 500
rect -1168 -488 -1162 488
rect -1128 -488 -1122 488
rect -1168 -500 -1122 -488
rect -710 488 -664 500
rect -710 -488 -704 488
rect -670 -488 -664 488
rect -710 -500 -664 -488
rect -252 488 -206 500
rect -252 -488 -246 488
rect -212 -488 -206 488
rect -252 -500 -206 -488
rect 206 488 252 500
rect 206 -488 212 488
rect 246 -488 252 488
rect 206 -500 252 -488
rect 664 488 710 500
rect 664 -488 670 488
rect 704 -488 710 488
rect 664 -500 710 -488
rect 1122 488 1168 500
rect 1122 -488 1128 488
rect 1162 -488 1168 488
rect 1122 -500 1168 -488
rect 1580 488 1626 500
rect 1580 -488 1586 488
rect 1620 -488 1626 488
rect 1580 -500 1626 -488
rect 2038 488 2084 500
rect 2038 -488 2044 488
rect 2078 -488 2084 488
rect 2038 -500 2084 -488
rect -2028 -547 -1636 -541
rect -2028 -581 -2016 -547
rect -1648 -581 -1636 -547
rect -2028 -587 -1636 -581
rect -1570 -547 -1178 -541
rect -1570 -581 -1558 -547
rect -1190 -581 -1178 -547
rect -1570 -587 -1178 -581
rect -1112 -547 -720 -541
rect -1112 -581 -1100 -547
rect -732 -581 -720 -547
rect -1112 -587 -720 -581
rect -654 -547 -262 -541
rect -654 -581 -642 -547
rect -274 -581 -262 -547
rect -654 -587 -262 -581
rect -196 -547 196 -541
rect -196 -581 -184 -547
rect 184 -581 196 -547
rect -196 -587 196 -581
rect 262 -547 654 -541
rect 262 -581 274 -547
rect 642 -581 654 -547
rect 262 -587 654 -581
rect 720 -547 1112 -541
rect 720 -581 732 -547
rect 1100 -581 1112 -547
rect 720 -587 1112 -581
rect 1178 -547 1570 -541
rect 1178 -581 1190 -547
rect 1558 -581 1570 -547
rect 1178 -587 1570 -581
rect 1636 -547 2028 -541
rect 1636 -581 1648 -547
rect 2016 -581 2028 -547
rect 1636 -587 2028 -581
<< properties >>
string FIXED_BBOX -2195 -702 2195 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 2 m 1 nf 9 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
