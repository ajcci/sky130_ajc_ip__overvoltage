magic
tech sky130A
magscale 1 2
timestamp 1711685078
<< error_p >>
rect 20177 -5347 20205 -5345
rect 20177 -5365 20219 -5347
rect 20157 -5369 20225 -5365
rect 20157 -5389 20215 -5369
rect 20219 -5389 20225 -5369
rect 20157 -5393 20225 -5389
rect 20177 -5405 20219 -5393
rect 20177 -5413 20205 -5405
<< error_s >>
rect 19966 -1772 20028 -1766
rect 19966 -1806 19982 -1772
rect 19966 -1812 20028 -1806
rect 19970 -1966 20028 -1960
rect 19970 -2000 19982 -1966
rect 19970 -2006 20028 -2000
<< dnwell >>
rect 8363 -9837 36013 3064
<< nwell >>
rect 8283 2858 36093 3144
rect 8283 -9631 8569 2858
rect 35807 -9631 36093 2858
rect 8283 -9917 36093 -9631
<< pwell >>
rect 4522 -3169 6500 -1640
rect 16688 -5933 24802 523
<< nsubdiff >>
rect 8320 3087 36056 3107
rect 8320 3053 8400 3087
rect 35976 3053 36056 3087
rect 8320 3033 36056 3053
rect 8320 3027 8394 3033
rect 8320 -9800 8340 3027
rect 8374 -9800 8394 3027
rect 35982 3027 36056 3033
rect 8320 -9806 8394 -9800
rect 35982 -9800 36002 3027
rect 36036 -9800 36056 3027
rect 35982 -9806 36056 -9800
rect 8320 -9826 36056 -9806
rect 8320 -9860 8400 -9826
rect 35976 -9860 36056 -9826
rect 8320 -9880 36056 -9860
<< mvpsubdiff >>
rect 5484 -2434 5665 -2401
rect 5484 -2468 5541 -2434
rect 5605 -2468 5665 -2434
rect 5484 -2492 5665 -2468
rect 20181 -5369 20219 -5347
rect 20201 -5389 20219 -5369
rect 20181 -5405 20219 -5389
<< nsubdiffcont >>
rect 8400 3053 35976 3087
rect 8340 -9800 8374 3027
rect 36002 -9800 36036 3027
rect 8400 -9860 35976 -9826
<< mvpsubdiffcont >>
rect 5541 -2468 5605 -2434
rect 20181 -5389 20201 -5369
<< locali >>
rect 8340 3053 8400 3087
rect 35976 3053 36036 3087
rect 8340 3027 8374 3053
rect 5516 -2434 5627 -2420
rect 5516 -2468 5541 -2434
rect 5605 -2468 5627 -2434
rect 5516 -2480 5627 -2468
rect 5547 -2520 5584 -2480
rect 36002 3027 36036 3053
rect 20231 -5359 20265 -5297
rect 19839 -5369 20265 -5359
rect 19839 -5389 20181 -5369
rect 20201 -5389 20265 -5369
rect 19839 -5393 20265 -5389
rect 8340 -9826 8374 -9800
rect 36002 -9826 36036 -9800
rect 8340 -9860 8400 -9826
rect 35976 -9860 36036 -9826
<< viali >>
rect 8340 -2485 8374 -2423
<< metal1 >>
rect 19966 -1812 19970 -1766
rect 19932 -1844 19978 -1840
rect 20020 -1844 20066 -1840
rect 8329 -2423 8385 -2409
rect 8329 -2485 8340 -2423
rect 8374 -2485 8385 -2423
rect 8329 -2497 8385 -2485
use sky130_fd_pr__nfet_01v8_7XH9KL  sky130_fd_pr__nfet_01v8_7XH9KL_0
timestamp 1711685078
transform 1 0 19999 0 1 -1886
box -73 -130 73 130
<< labels >>
rlabel metal1 8329 -2444 8329 -2444 1 avdd
port 0 n
rlabel locali 5547 -2520 5547 -2520 1 avss
rlabel locali 20248 -5338 20248 -5338 1 vt
rlabel metal1 19966 -1766 19966 -1766 1 g
rlabel metal1 19932 -1840 19932 -1840 1 d
rlabel metal1 20066 -1840 20066 -1840 1 s
<< end >>
