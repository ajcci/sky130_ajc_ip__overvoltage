magic
tech sky130A
magscale 1 2
timestamp 1711568248
<< pwell >>
rect -8489 -753 8489 753
<< mvnmos >>
rect -8261 411 -6661 495
rect -6603 411 -5003 495
rect -4945 411 -3345 495
rect -3287 411 -1687 495
rect -1629 411 -29 495
rect 29 411 1629 495
rect 1687 411 3287 495
rect 3345 411 4945 495
rect 5003 411 6603 495
rect 6661 411 8261 495
rect -8261 109 -6661 193
rect -6603 109 -5003 193
rect -4945 109 -3345 193
rect -3287 109 -1687 193
rect -1629 109 -29 193
rect 29 109 1629 193
rect 1687 109 3287 193
rect 3345 109 4945 193
rect 5003 109 6603 193
rect 6661 109 8261 193
rect -8261 -193 -6661 -109
rect -6603 -193 -5003 -109
rect -4945 -193 -3345 -109
rect -3287 -193 -1687 -109
rect -1629 -193 -29 -109
rect 29 -193 1629 -109
rect 1687 -193 3287 -109
rect 3345 -193 4945 -109
rect 5003 -193 6603 -109
rect 6661 -193 8261 -109
rect -8261 -495 -6661 -411
rect -6603 -495 -5003 -411
rect -4945 -495 -3345 -411
rect -3287 -495 -1687 -411
rect -1629 -495 -29 -411
rect 29 -495 1629 -411
rect 1687 -495 3287 -411
rect 3345 -495 4945 -411
rect 5003 -495 6603 -411
rect 6661 -495 8261 -411
<< mvndiff >>
rect -8319 483 -8261 495
rect -8319 423 -8307 483
rect -8273 423 -8261 483
rect -8319 411 -8261 423
rect -6661 483 -6603 495
rect -6661 423 -6649 483
rect -6615 423 -6603 483
rect -6661 411 -6603 423
rect -5003 483 -4945 495
rect -5003 423 -4991 483
rect -4957 423 -4945 483
rect -5003 411 -4945 423
rect -3345 483 -3287 495
rect -3345 423 -3333 483
rect -3299 423 -3287 483
rect -3345 411 -3287 423
rect -1687 483 -1629 495
rect -1687 423 -1675 483
rect -1641 423 -1629 483
rect -1687 411 -1629 423
rect -29 483 29 495
rect -29 423 -17 483
rect 17 423 29 483
rect -29 411 29 423
rect 1629 483 1687 495
rect 1629 423 1641 483
rect 1675 423 1687 483
rect 1629 411 1687 423
rect 3287 483 3345 495
rect 3287 423 3299 483
rect 3333 423 3345 483
rect 3287 411 3345 423
rect 4945 483 5003 495
rect 4945 423 4957 483
rect 4991 423 5003 483
rect 4945 411 5003 423
rect 6603 483 6661 495
rect 6603 423 6615 483
rect 6649 423 6661 483
rect 6603 411 6661 423
rect 8261 483 8319 495
rect 8261 423 8273 483
rect 8307 423 8319 483
rect 8261 411 8319 423
rect -8319 181 -8261 193
rect -8319 121 -8307 181
rect -8273 121 -8261 181
rect -8319 109 -8261 121
rect -6661 181 -6603 193
rect -6661 121 -6649 181
rect -6615 121 -6603 181
rect -6661 109 -6603 121
rect -5003 181 -4945 193
rect -5003 121 -4991 181
rect -4957 121 -4945 181
rect -5003 109 -4945 121
rect -3345 181 -3287 193
rect -3345 121 -3333 181
rect -3299 121 -3287 181
rect -3345 109 -3287 121
rect -1687 181 -1629 193
rect -1687 121 -1675 181
rect -1641 121 -1629 181
rect -1687 109 -1629 121
rect -29 181 29 193
rect -29 121 -17 181
rect 17 121 29 181
rect -29 109 29 121
rect 1629 181 1687 193
rect 1629 121 1641 181
rect 1675 121 1687 181
rect 1629 109 1687 121
rect 3287 181 3345 193
rect 3287 121 3299 181
rect 3333 121 3345 181
rect 3287 109 3345 121
rect 4945 181 5003 193
rect 4945 121 4957 181
rect 4991 121 5003 181
rect 4945 109 5003 121
rect 6603 181 6661 193
rect 6603 121 6615 181
rect 6649 121 6661 181
rect 6603 109 6661 121
rect 8261 181 8319 193
rect 8261 121 8273 181
rect 8307 121 8319 181
rect 8261 109 8319 121
rect -8319 -121 -8261 -109
rect -8319 -181 -8307 -121
rect -8273 -181 -8261 -121
rect -8319 -193 -8261 -181
rect -6661 -121 -6603 -109
rect -6661 -181 -6649 -121
rect -6615 -181 -6603 -121
rect -6661 -193 -6603 -181
rect -5003 -121 -4945 -109
rect -5003 -181 -4991 -121
rect -4957 -181 -4945 -121
rect -5003 -193 -4945 -181
rect -3345 -121 -3287 -109
rect -3345 -181 -3333 -121
rect -3299 -181 -3287 -121
rect -3345 -193 -3287 -181
rect -1687 -121 -1629 -109
rect -1687 -181 -1675 -121
rect -1641 -181 -1629 -121
rect -1687 -193 -1629 -181
rect -29 -121 29 -109
rect -29 -181 -17 -121
rect 17 -181 29 -121
rect -29 -193 29 -181
rect 1629 -121 1687 -109
rect 1629 -181 1641 -121
rect 1675 -181 1687 -121
rect 1629 -193 1687 -181
rect 3287 -121 3345 -109
rect 3287 -181 3299 -121
rect 3333 -181 3345 -121
rect 3287 -193 3345 -181
rect 4945 -121 5003 -109
rect 4945 -181 4957 -121
rect 4991 -181 5003 -121
rect 4945 -193 5003 -181
rect 6603 -121 6661 -109
rect 6603 -181 6615 -121
rect 6649 -181 6661 -121
rect 6603 -193 6661 -181
rect 8261 -121 8319 -109
rect 8261 -181 8273 -121
rect 8307 -181 8319 -121
rect 8261 -193 8319 -181
rect -8319 -423 -8261 -411
rect -8319 -483 -8307 -423
rect -8273 -483 -8261 -423
rect -8319 -495 -8261 -483
rect -6661 -423 -6603 -411
rect -6661 -483 -6649 -423
rect -6615 -483 -6603 -423
rect -6661 -495 -6603 -483
rect -5003 -423 -4945 -411
rect -5003 -483 -4991 -423
rect -4957 -483 -4945 -423
rect -5003 -495 -4945 -483
rect -3345 -423 -3287 -411
rect -3345 -483 -3333 -423
rect -3299 -483 -3287 -423
rect -3345 -495 -3287 -483
rect -1687 -423 -1629 -411
rect -1687 -483 -1675 -423
rect -1641 -483 -1629 -423
rect -1687 -495 -1629 -483
rect -29 -423 29 -411
rect -29 -483 -17 -423
rect 17 -483 29 -423
rect -29 -495 29 -483
rect 1629 -423 1687 -411
rect 1629 -483 1641 -423
rect 1675 -483 1687 -423
rect 1629 -495 1687 -483
rect 3287 -423 3345 -411
rect 3287 -483 3299 -423
rect 3333 -483 3345 -423
rect 3287 -495 3345 -483
rect 4945 -423 5003 -411
rect 4945 -483 4957 -423
rect 4991 -483 5003 -423
rect 4945 -495 5003 -483
rect 6603 -423 6661 -411
rect 6603 -483 6615 -423
rect 6649 -483 6661 -423
rect 6603 -495 6661 -483
rect 8261 -423 8319 -411
rect 8261 -483 8273 -423
rect 8307 -483 8319 -423
rect 8261 -495 8319 -483
<< mvndiffc >>
rect -8307 423 -8273 483
rect -6649 423 -6615 483
rect -4991 423 -4957 483
rect -3333 423 -3299 483
rect -1675 423 -1641 483
rect -17 423 17 483
rect 1641 423 1675 483
rect 3299 423 3333 483
rect 4957 423 4991 483
rect 6615 423 6649 483
rect 8273 423 8307 483
rect -8307 121 -8273 181
rect -6649 121 -6615 181
rect -4991 121 -4957 181
rect -3333 121 -3299 181
rect -1675 121 -1641 181
rect -17 121 17 181
rect 1641 121 1675 181
rect 3299 121 3333 181
rect 4957 121 4991 181
rect 6615 121 6649 181
rect 8273 121 8307 181
rect -8307 -181 -8273 -121
rect -6649 -181 -6615 -121
rect -4991 -181 -4957 -121
rect -3333 -181 -3299 -121
rect -1675 -181 -1641 -121
rect -17 -181 17 -121
rect 1641 -181 1675 -121
rect 3299 -181 3333 -121
rect 4957 -181 4991 -121
rect 6615 -181 6649 -121
rect 8273 -181 8307 -121
rect -8307 -483 -8273 -423
rect -6649 -483 -6615 -423
rect -4991 -483 -4957 -423
rect -3333 -483 -3299 -423
rect -1675 -483 -1641 -423
rect -17 -483 17 -423
rect 1641 -483 1675 -423
rect 3299 -483 3333 -423
rect 4957 -483 4991 -423
rect 6615 -483 6649 -423
rect 8273 -483 8307 -423
<< mvpsubdiff >>
rect -8453 705 8453 717
rect -8453 671 -8345 705
rect 8345 671 8453 705
rect -8453 659 8453 671
rect -8453 609 -8395 659
rect -8453 -609 -8441 609
rect -8407 -609 -8395 609
rect 8395 609 8453 659
rect -8453 -659 -8395 -609
rect 8395 -609 8407 609
rect 8441 -609 8453 609
rect 8395 -659 8453 -609
rect -8453 -671 8453 -659
rect -8453 -705 -8345 -671
rect 8345 -705 8453 -671
rect -8453 -717 8453 -705
<< mvpsubdiffcont >>
rect -8345 671 8345 705
rect -8441 -609 -8407 609
rect 8407 -609 8441 609
rect -8345 -705 8345 -671
<< poly >>
rect -8261 567 -6661 583
rect -8261 533 -8245 567
rect -6677 533 -6661 567
rect -8261 495 -6661 533
rect -6603 567 -5003 583
rect -6603 533 -6587 567
rect -5019 533 -5003 567
rect -6603 495 -5003 533
rect -4945 567 -3345 583
rect -4945 533 -4929 567
rect -3361 533 -3345 567
rect -4945 495 -3345 533
rect -3287 567 -1687 583
rect -3287 533 -3271 567
rect -1703 533 -1687 567
rect -3287 495 -1687 533
rect -1629 567 -29 583
rect -1629 533 -1613 567
rect -45 533 -29 567
rect -1629 495 -29 533
rect 29 567 1629 583
rect 29 533 45 567
rect 1613 533 1629 567
rect 29 495 1629 533
rect 1687 567 3287 583
rect 1687 533 1703 567
rect 3271 533 3287 567
rect 1687 495 3287 533
rect 3345 567 4945 583
rect 3345 533 3361 567
rect 4929 533 4945 567
rect 3345 495 4945 533
rect 5003 567 6603 583
rect 5003 533 5019 567
rect 6587 533 6603 567
rect 5003 495 6603 533
rect 6661 567 8261 583
rect 6661 533 6677 567
rect 8245 533 8261 567
rect 6661 495 8261 533
rect -8261 373 -6661 411
rect -8261 339 -8245 373
rect -6677 339 -6661 373
rect -8261 323 -6661 339
rect -6603 373 -5003 411
rect -6603 339 -6587 373
rect -5019 339 -5003 373
rect -6603 323 -5003 339
rect -4945 373 -3345 411
rect -4945 339 -4929 373
rect -3361 339 -3345 373
rect -4945 323 -3345 339
rect -3287 373 -1687 411
rect -3287 339 -3271 373
rect -1703 339 -1687 373
rect -3287 323 -1687 339
rect -1629 373 -29 411
rect -1629 339 -1613 373
rect -45 339 -29 373
rect -1629 323 -29 339
rect 29 373 1629 411
rect 29 339 45 373
rect 1613 339 1629 373
rect 29 323 1629 339
rect 1687 373 3287 411
rect 1687 339 1703 373
rect 3271 339 3287 373
rect 1687 323 3287 339
rect 3345 373 4945 411
rect 3345 339 3361 373
rect 4929 339 4945 373
rect 3345 323 4945 339
rect 5003 373 6603 411
rect 5003 339 5019 373
rect 6587 339 6603 373
rect 5003 323 6603 339
rect 6661 373 8261 411
rect 6661 339 6677 373
rect 8245 339 8261 373
rect 6661 323 8261 339
rect -8261 265 -6661 281
rect -8261 231 -8245 265
rect -6677 231 -6661 265
rect -8261 193 -6661 231
rect -6603 265 -5003 281
rect -6603 231 -6587 265
rect -5019 231 -5003 265
rect -6603 193 -5003 231
rect -4945 265 -3345 281
rect -4945 231 -4929 265
rect -3361 231 -3345 265
rect -4945 193 -3345 231
rect -3287 265 -1687 281
rect -3287 231 -3271 265
rect -1703 231 -1687 265
rect -3287 193 -1687 231
rect -1629 265 -29 281
rect -1629 231 -1613 265
rect -45 231 -29 265
rect -1629 193 -29 231
rect 29 265 1629 281
rect 29 231 45 265
rect 1613 231 1629 265
rect 29 193 1629 231
rect 1687 265 3287 281
rect 1687 231 1703 265
rect 3271 231 3287 265
rect 1687 193 3287 231
rect 3345 265 4945 281
rect 3345 231 3361 265
rect 4929 231 4945 265
rect 3345 193 4945 231
rect 5003 265 6603 281
rect 5003 231 5019 265
rect 6587 231 6603 265
rect 5003 193 6603 231
rect 6661 265 8261 281
rect 6661 231 6677 265
rect 8245 231 8261 265
rect 6661 193 8261 231
rect -8261 71 -6661 109
rect -8261 37 -8245 71
rect -6677 37 -6661 71
rect -8261 21 -6661 37
rect -6603 71 -5003 109
rect -6603 37 -6587 71
rect -5019 37 -5003 71
rect -6603 21 -5003 37
rect -4945 71 -3345 109
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -4945 21 -3345 37
rect -3287 71 -1687 109
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -3287 21 -1687 37
rect -1629 71 -29 109
rect -1629 37 -1613 71
rect -45 37 -29 71
rect -1629 21 -29 37
rect 29 71 1629 109
rect 29 37 45 71
rect 1613 37 1629 71
rect 29 21 1629 37
rect 1687 71 3287 109
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 1687 21 3287 37
rect 3345 71 4945 109
rect 3345 37 3361 71
rect 4929 37 4945 71
rect 3345 21 4945 37
rect 5003 71 6603 109
rect 5003 37 5019 71
rect 6587 37 6603 71
rect 5003 21 6603 37
rect 6661 71 8261 109
rect 6661 37 6677 71
rect 8245 37 8261 71
rect 6661 21 8261 37
rect -8261 -37 -6661 -21
rect -8261 -71 -8245 -37
rect -6677 -71 -6661 -37
rect -8261 -109 -6661 -71
rect -6603 -37 -5003 -21
rect -6603 -71 -6587 -37
rect -5019 -71 -5003 -37
rect -6603 -109 -5003 -71
rect -4945 -37 -3345 -21
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -4945 -109 -3345 -71
rect -3287 -37 -1687 -21
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -3287 -109 -1687 -71
rect -1629 -37 -29 -21
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect -1629 -109 -29 -71
rect 29 -37 1629 -21
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 29 -109 1629 -71
rect 1687 -37 3287 -21
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 1687 -109 3287 -71
rect 3345 -37 4945 -21
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect 3345 -109 4945 -71
rect 5003 -37 6603 -21
rect 5003 -71 5019 -37
rect 6587 -71 6603 -37
rect 5003 -109 6603 -71
rect 6661 -37 8261 -21
rect 6661 -71 6677 -37
rect 8245 -71 8261 -37
rect 6661 -109 8261 -71
rect -8261 -231 -6661 -193
rect -8261 -265 -8245 -231
rect -6677 -265 -6661 -231
rect -8261 -281 -6661 -265
rect -6603 -231 -5003 -193
rect -6603 -265 -6587 -231
rect -5019 -265 -5003 -231
rect -6603 -281 -5003 -265
rect -4945 -231 -3345 -193
rect -4945 -265 -4929 -231
rect -3361 -265 -3345 -231
rect -4945 -281 -3345 -265
rect -3287 -231 -1687 -193
rect -3287 -265 -3271 -231
rect -1703 -265 -1687 -231
rect -3287 -281 -1687 -265
rect -1629 -231 -29 -193
rect -1629 -265 -1613 -231
rect -45 -265 -29 -231
rect -1629 -281 -29 -265
rect 29 -231 1629 -193
rect 29 -265 45 -231
rect 1613 -265 1629 -231
rect 29 -281 1629 -265
rect 1687 -231 3287 -193
rect 1687 -265 1703 -231
rect 3271 -265 3287 -231
rect 1687 -281 3287 -265
rect 3345 -231 4945 -193
rect 3345 -265 3361 -231
rect 4929 -265 4945 -231
rect 3345 -281 4945 -265
rect 5003 -231 6603 -193
rect 5003 -265 5019 -231
rect 6587 -265 6603 -231
rect 5003 -281 6603 -265
rect 6661 -231 8261 -193
rect 6661 -265 6677 -231
rect 8245 -265 8261 -231
rect 6661 -281 8261 -265
rect -8261 -339 -6661 -323
rect -8261 -373 -8245 -339
rect -6677 -373 -6661 -339
rect -8261 -411 -6661 -373
rect -6603 -339 -5003 -323
rect -6603 -373 -6587 -339
rect -5019 -373 -5003 -339
rect -6603 -411 -5003 -373
rect -4945 -339 -3345 -323
rect -4945 -373 -4929 -339
rect -3361 -373 -3345 -339
rect -4945 -411 -3345 -373
rect -3287 -339 -1687 -323
rect -3287 -373 -3271 -339
rect -1703 -373 -1687 -339
rect -3287 -411 -1687 -373
rect -1629 -339 -29 -323
rect -1629 -373 -1613 -339
rect -45 -373 -29 -339
rect -1629 -411 -29 -373
rect 29 -339 1629 -323
rect 29 -373 45 -339
rect 1613 -373 1629 -339
rect 29 -411 1629 -373
rect 1687 -339 3287 -323
rect 1687 -373 1703 -339
rect 3271 -373 3287 -339
rect 1687 -411 3287 -373
rect 3345 -339 4945 -323
rect 3345 -373 3361 -339
rect 4929 -373 4945 -339
rect 3345 -411 4945 -373
rect 5003 -339 6603 -323
rect 5003 -373 5019 -339
rect 6587 -373 6603 -339
rect 5003 -411 6603 -373
rect 6661 -339 8261 -323
rect 6661 -373 6677 -339
rect 8245 -373 8261 -339
rect 6661 -411 8261 -373
rect -8261 -533 -6661 -495
rect -8261 -567 -8245 -533
rect -6677 -567 -6661 -533
rect -8261 -583 -6661 -567
rect -6603 -533 -5003 -495
rect -6603 -567 -6587 -533
rect -5019 -567 -5003 -533
rect -6603 -583 -5003 -567
rect -4945 -533 -3345 -495
rect -4945 -567 -4929 -533
rect -3361 -567 -3345 -533
rect -4945 -583 -3345 -567
rect -3287 -533 -1687 -495
rect -3287 -567 -3271 -533
rect -1703 -567 -1687 -533
rect -3287 -583 -1687 -567
rect -1629 -533 -29 -495
rect -1629 -567 -1613 -533
rect -45 -567 -29 -533
rect -1629 -583 -29 -567
rect 29 -533 1629 -495
rect 29 -567 45 -533
rect 1613 -567 1629 -533
rect 29 -583 1629 -567
rect 1687 -533 3287 -495
rect 1687 -567 1703 -533
rect 3271 -567 3287 -533
rect 1687 -583 3287 -567
rect 3345 -533 4945 -495
rect 3345 -567 3361 -533
rect 4929 -567 4945 -533
rect 3345 -583 4945 -567
rect 5003 -533 6603 -495
rect 5003 -567 5019 -533
rect 6587 -567 6603 -533
rect 5003 -583 6603 -567
rect 6661 -533 8261 -495
rect 6661 -567 6677 -533
rect 8245 -567 8261 -533
rect 6661 -583 8261 -567
<< polycont >>
rect -8245 533 -6677 567
rect -6587 533 -5019 567
rect -4929 533 -3361 567
rect -3271 533 -1703 567
rect -1613 533 -45 567
rect 45 533 1613 567
rect 1703 533 3271 567
rect 3361 533 4929 567
rect 5019 533 6587 567
rect 6677 533 8245 567
rect -8245 339 -6677 373
rect -6587 339 -5019 373
rect -4929 339 -3361 373
rect -3271 339 -1703 373
rect -1613 339 -45 373
rect 45 339 1613 373
rect 1703 339 3271 373
rect 3361 339 4929 373
rect 5019 339 6587 373
rect 6677 339 8245 373
rect -8245 231 -6677 265
rect -6587 231 -5019 265
rect -4929 231 -3361 265
rect -3271 231 -1703 265
rect -1613 231 -45 265
rect 45 231 1613 265
rect 1703 231 3271 265
rect 3361 231 4929 265
rect 5019 231 6587 265
rect 6677 231 8245 265
rect -8245 37 -6677 71
rect -6587 37 -5019 71
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect 5019 37 6587 71
rect 6677 37 8245 71
rect -8245 -71 -6677 -37
rect -6587 -71 -5019 -37
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
rect 5019 -71 6587 -37
rect 6677 -71 8245 -37
rect -8245 -265 -6677 -231
rect -6587 -265 -5019 -231
rect -4929 -265 -3361 -231
rect -3271 -265 -1703 -231
rect -1613 -265 -45 -231
rect 45 -265 1613 -231
rect 1703 -265 3271 -231
rect 3361 -265 4929 -231
rect 5019 -265 6587 -231
rect 6677 -265 8245 -231
rect -8245 -373 -6677 -339
rect -6587 -373 -5019 -339
rect -4929 -373 -3361 -339
rect -3271 -373 -1703 -339
rect -1613 -373 -45 -339
rect 45 -373 1613 -339
rect 1703 -373 3271 -339
rect 3361 -373 4929 -339
rect 5019 -373 6587 -339
rect 6677 -373 8245 -339
rect -8245 -567 -6677 -533
rect -6587 -567 -5019 -533
rect -4929 -567 -3361 -533
rect -3271 -567 -1703 -533
rect -1613 -567 -45 -533
rect 45 -567 1613 -533
rect 1703 -567 3271 -533
rect 3361 -567 4929 -533
rect 5019 -567 6587 -533
rect 6677 -567 8245 -533
<< locali >>
rect -8441 671 -8345 705
rect 8345 671 8441 705
rect -8441 609 -8407 671
rect 8407 609 8441 671
rect -8261 533 -8245 567
rect -6677 533 -6661 567
rect -6603 533 -6587 567
rect -5019 533 -5003 567
rect -4945 533 -4929 567
rect -3361 533 -3345 567
rect -3287 533 -3271 567
rect -1703 533 -1687 567
rect -1629 533 -1613 567
rect -45 533 -29 567
rect 29 533 45 567
rect 1613 533 1629 567
rect 1687 533 1703 567
rect 3271 533 3287 567
rect 3345 533 3361 567
rect 4929 533 4945 567
rect 5003 533 5019 567
rect 6587 533 6603 567
rect 6661 533 6677 567
rect 8245 533 8261 567
rect -8307 483 -8273 499
rect -8307 407 -8273 423
rect -6649 483 -6615 499
rect -6649 407 -6615 423
rect -4991 483 -4957 499
rect -4991 407 -4957 423
rect -3333 483 -3299 499
rect -3333 407 -3299 423
rect -1675 483 -1641 499
rect -1675 407 -1641 423
rect -17 483 17 499
rect -17 407 17 423
rect 1641 483 1675 499
rect 1641 407 1675 423
rect 3299 483 3333 499
rect 3299 407 3333 423
rect 4957 483 4991 499
rect 4957 407 4991 423
rect 6615 483 6649 499
rect 6615 407 6649 423
rect 8273 483 8307 499
rect 8273 407 8307 423
rect -8261 339 -8245 373
rect -6677 339 -6661 373
rect -6603 339 -6587 373
rect -5019 339 -5003 373
rect -4945 339 -4929 373
rect -3361 339 -3345 373
rect -3287 339 -3271 373
rect -1703 339 -1687 373
rect -1629 339 -1613 373
rect -45 339 -29 373
rect 29 339 45 373
rect 1613 339 1629 373
rect 1687 339 1703 373
rect 3271 339 3287 373
rect 3345 339 3361 373
rect 4929 339 4945 373
rect 5003 339 5019 373
rect 6587 339 6603 373
rect 6661 339 6677 373
rect 8245 339 8261 373
rect -8261 231 -8245 265
rect -6677 231 -6661 265
rect -6603 231 -6587 265
rect -5019 231 -5003 265
rect -4945 231 -4929 265
rect -3361 231 -3345 265
rect -3287 231 -3271 265
rect -1703 231 -1687 265
rect -1629 231 -1613 265
rect -45 231 -29 265
rect 29 231 45 265
rect 1613 231 1629 265
rect 1687 231 1703 265
rect 3271 231 3287 265
rect 3345 231 3361 265
rect 4929 231 4945 265
rect 5003 231 5019 265
rect 6587 231 6603 265
rect 6661 231 6677 265
rect 8245 231 8261 265
rect -8307 181 -8273 197
rect -8307 105 -8273 121
rect -6649 181 -6615 197
rect -6649 105 -6615 121
rect -4991 181 -4957 197
rect -4991 105 -4957 121
rect -3333 181 -3299 197
rect -3333 105 -3299 121
rect -1675 181 -1641 197
rect -1675 105 -1641 121
rect -17 181 17 197
rect -17 105 17 121
rect 1641 181 1675 197
rect 1641 105 1675 121
rect 3299 181 3333 197
rect 3299 105 3333 121
rect 4957 181 4991 197
rect 4957 105 4991 121
rect 6615 181 6649 197
rect 6615 105 6649 121
rect 8273 181 8307 197
rect 8273 105 8307 121
rect -8261 37 -8245 71
rect -6677 37 -6661 71
rect -6603 37 -6587 71
rect -5019 37 -5003 71
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -1629 37 -1613 71
rect -45 37 -29 71
rect 29 37 45 71
rect 1613 37 1629 71
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 3345 37 3361 71
rect 4929 37 4945 71
rect 5003 37 5019 71
rect 6587 37 6603 71
rect 6661 37 6677 71
rect 8245 37 8261 71
rect -8261 -71 -8245 -37
rect -6677 -71 -6661 -37
rect -6603 -71 -6587 -37
rect -5019 -71 -5003 -37
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect 5003 -71 5019 -37
rect 6587 -71 6603 -37
rect 6661 -71 6677 -37
rect 8245 -71 8261 -37
rect -8307 -121 -8273 -105
rect -8307 -197 -8273 -181
rect -6649 -121 -6615 -105
rect -6649 -197 -6615 -181
rect -4991 -121 -4957 -105
rect -4991 -197 -4957 -181
rect -3333 -121 -3299 -105
rect -3333 -197 -3299 -181
rect -1675 -121 -1641 -105
rect -1675 -197 -1641 -181
rect -17 -121 17 -105
rect -17 -197 17 -181
rect 1641 -121 1675 -105
rect 1641 -197 1675 -181
rect 3299 -121 3333 -105
rect 3299 -197 3333 -181
rect 4957 -121 4991 -105
rect 4957 -197 4991 -181
rect 6615 -121 6649 -105
rect 6615 -197 6649 -181
rect 8273 -121 8307 -105
rect 8273 -197 8307 -181
rect -8261 -265 -8245 -231
rect -6677 -265 -6661 -231
rect -6603 -265 -6587 -231
rect -5019 -265 -5003 -231
rect -4945 -265 -4929 -231
rect -3361 -265 -3345 -231
rect -3287 -265 -3271 -231
rect -1703 -265 -1687 -231
rect -1629 -265 -1613 -231
rect -45 -265 -29 -231
rect 29 -265 45 -231
rect 1613 -265 1629 -231
rect 1687 -265 1703 -231
rect 3271 -265 3287 -231
rect 3345 -265 3361 -231
rect 4929 -265 4945 -231
rect 5003 -265 5019 -231
rect 6587 -265 6603 -231
rect 6661 -265 6677 -231
rect 8245 -265 8261 -231
rect -8261 -373 -8245 -339
rect -6677 -373 -6661 -339
rect -6603 -373 -6587 -339
rect -5019 -373 -5003 -339
rect -4945 -373 -4929 -339
rect -3361 -373 -3345 -339
rect -3287 -373 -3271 -339
rect -1703 -373 -1687 -339
rect -1629 -373 -1613 -339
rect -45 -373 -29 -339
rect 29 -373 45 -339
rect 1613 -373 1629 -339
rect 1687 -373 1703 -339
rect 3271 -373 3287 -339
rect 3345 -373 3361 -339
rect 4929 -373 4945 -339
rect 5003 -373 5019 -339
rect 6587 -373 6603 -339
rect 6661 -373 6677 -339
rect 8245 -373 8261 -339
rect -8307 -423 -8273 -407
rect -8307 -499 -8273 -483
rect -6649 -423 -6615 -407
rect -6649 -499 -6615 -483
rect -4991 -423 -4957 -407
rect -4991 -499 -4957 -483
rect -3333 -423 -3299 -407
rect -3333 -499 -3299 -483
rect -1675 -423 -1641 -407
rect -1675 -499 -1641 -483
rect -17 -423 17 -407
rect -17 -499 17 -483
rect 1641 -423 1675 -407
rect 1641 -499 1675 -483
rect 3299 -423 3333 -407
rect 3299 -499 3333 -483
rect 4957 -423 4991 -407
rect 4957 -499 4991 -483
rect 6615 -423 6649 -407
rect 6615 -499 6649 -483
rect 8273 -423 8307 -407
rect 8273 -499 8307 -483
rect -8261 -567 -8245 -533
rect -6677 -567 -6661 -533
rect -6603 -567 -6587 -533
rect -5019 -567 -5003 -533
rect -4945 -567 -4929 -533
rect -3361 -567 -3345 -533
rect -3287 -567 -3271 -533
rect -1703 -567 -1687 -533
rect -1629 -567 -1613 -533
rect -45 -567 -29 -533
rect 29 -567 45 -533
rect 1613 -567 1629 -533
rect 1687 -567 1703 -533
rect 3271 -567 3287 -533
rect 3345 -567 3361 -533
rect 4929 -567 4945 -533
rect 5003 -567 5019 -533
rect 6587 -567 6603 -533
rect 6661 -567 6677 -533
rect 8245 -567 8261 -533
rect -8441 -671 -8407 -609
rect 8407 -671 8441 -609
rect -8441 -705 -8345 -671
rect 8345 -705 8441 -671
<< viali >>
rect -8245 533 -6677 567
rect -6587 533 -5019 567
rect -4929 533 -3361 567
rect -3271 533 -1703 567
rect -1613 533 -45 567
rect 45 533 1613 567
rect 1703 533 3271 567
rect 3361 533 4929 567
rect 5019 533 6587 567
rect 6677 533 8245 567
rect -8307 423 -8273 483
rect -6649 423 -6615 483
rect -4991 423 -4957 483
rect -3333 423 -3299 483
rect -1675 423 -1641 483
rect -17 423 17 483
rect 1641 423 1675 483
rect 3299 423 3333 483
rect 4957 423 4991 483
rect 6615 423 6649 483
rect 8273 423 8307 483
rect -8245 339 -6677 373
rect -6587 339 -5019 373
rect -4929 339 -3361 373
rect -3271 339 -1703 373
rect -1613 339 -45 373
rect 45 339 1613 373
rect 1703 339 3271 373
rect 3361 339 4929 373
rect 5019 339 6587 373
rect 6677 339 8245 373
rect -8245 231 -6677 265
rect -6587 231 -5019 265
rect -4929 231 -3361 265
rect -3271 231 -1703 265
rect -1613 231 -45 265
rect 45 231 1613 265
rect 1703 231 3271 265
rect 3361 231 4929 265
rect 5019 231 6587 265
rect 6677 231 8245 265
rect -8307 121 -8273 181
rect -6649 121 -6615 181
rect -4991 121 -4957 181
rect -3333 121 -3299 181
rect -1675 121 -1641 181
rect -17 121 17 181
rect 1641 121 1675 181
rect 3299 121 3333 181
rect 4957 121 4991 181
rect 6615 121 6649 181
rect 8273 121 8307 181
rect -8245 37 -6677 71
rect -6587 37 -5019 71
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect 5019 37 6587 71
rect 6677 37 8245 71
rect -8245 -71 -6677 -37
rect -6587 -71 -5019 -37
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
rect 5019 -71 6587 -37
rect 6677 -71 8245 -37
rect -8307 -181 -8273 -121
rect -6649 -181 -6615 -121
rect -4991 -181 -4957 -121
rect -3333 -181 -3299 -121
rect -1675 -181 -1641 -121
rect -17 -181 17 -121
rect 1641 -181 1675 -121
rect 3299 -181 3333 -121
rect 4957 -181 4991 -121
rect 6615 -181 6649 -121
rect 8273 -181 8307 -121
rect -8245 -265 -6677 -231
rect -6587 -265 -5019 -231
rect -4929 -265 -3361 -231
rect -3271 -265 -1703 -231
rect -1613 -265 -45 -231
rect 45 -265 1613 -231
rect 1703 -265 3271 -231
rect 3361 -265 4929 -231
rect 5019 -265 6587 -231
rect 6677 -265 8245 -231
rect -8245 -373 -6677 -339
rect -6587 -373 -5019 -339
rect -4929 -373 -3361 -339
rect -3271 -373 -1703 -339
rect -1613 -373 -45 -339
rect 45 -373 1613 -339
rect 1703 -373 3271 -339
rect 3361 -373 4929 -339
rect 5019 -373 6587 -339
rect 6677 -373 8245 -339
rect -8307 -483 -8273 -423
rect -6649 -483 -6615 -423
rect -4991 -483 -4957 -423
rect -3333 -483 -3299 -423
rect -1675 -483 -1641 -423
rect -17 -483 17 -423
rect 1641 -483 1675 -423
rect 3299 -483 3333 -423
rect 4957 -483 4991 -423
rect 6615 -483 6649 -423
rect 8273 -483 8307 -423
rect -8245 -567 -6677 -533
rect -6587 -567 -5019 -533
rect -4929 -567 -3361 -533
rect -3271 -567 -1703 -533
rect -1613 -567 -45 -533
rect 45 -567 1613 -533
rect 1703 -567 3271 -533
rect 3361 -567 4929 -533
rect 5019 -567 6587 -533
rect 6677 -567 8245 -533
<< metal1 >>
rect -8257 567 -6665 573
rect -8257 533 -8245 567
rect -6677 533 -6665 567
rect -8257 527 -6665 533
rect -6599 567 -5007 573
rect -6599 533 -6587 567
rect -5019 533 -5007 567
rect -6599 527 -5007 533
rect -4941 567 -3349 573
rect -4941 533 -4929 567
rect -3361 533 -3349 567
rect -4941 527 -3349 533
rect -3283 567 -1691 573
rect -3283 533 -3271 567
rect -1703 533 -1691 567
rect -3283 527 -1691 533
rect -1625 567 -33 573
rect -1625 533 -1613 567
rect -45 533 -33 567
rect -1625 527 -33 533
rect 33 567 1625 573
rect 33 533 45 567
rect 1613 533 1625 567
rect 33 527 1625 533
rect 1691 567 3283 573
rect 1691 533 1703 567
rect 3271 533 3283 567
rect 1691 527 3283 533
rect 3349 567 4941 573
rect 3349 533 3361 567
rect 4929 533 4941 567
rect 3349 527 4941 533
rect 5007 567 6599 573
rect 5007 533 5019 567
rect 6587 533 6599 567
rect 5007 527 6599 533
rect 6665 567 8257 573
rect 6665 533 6677 567
rect 8245 533 8257 567
rect 6665 527 8257 533
rect -8313 483 -8267 495
rect -8313 423 -8307 483
rect -8273 423 -8267 483
rect -8313 411 -8267 423
rect -6655 483 -6609 495
rect -6655 423 -6649 483
rect -6615 423 -6609 483
rect -6655 411 -6609 423
rect -4997 483 -4951 495
rect -4997 423 -4991 483
rect -4957 423 -4951 483
rect -4997 411 -4951 423
rect -3339 483 -3293 495
rect -3339 423 -3333 483
rect -3299 423 -3293 483
rect -3339 411 -3293 423
rect -1681 483 -1635 495
rect -1681 423 -1675 483
rect -1641 423 -1635 483
rect -1681 411 -1635 423
rect -23 483 23 495
rect -23 423 -17 483
rect 17 423 23 483
rect -23 411 23 423
rect 1635 483 1681 495
rect 1635 423 1641 483
rect 1675 423 1681 483
rect 1635 411 1681 423
rect 3293 483 3339 495
rect 3293 423 3299 483
rect 3333 423 3339 483
rect 3293 411 3339 423
rect 4951 483 4997 495
rect 4951 423 4957 483
rect 4991 423 4997 483
rect 4951 411 4997 423
rect 6609 483 6655 495
rect 6609 423 6615 483
rect 6649 423 6655 483
rect 6609 411 6655 423
rect 8267 483 8313 495
rect 8267 423 8273 483
rect 8307 423 8313 483
rect 8267 411 8313 423
rect -8257 373 -6665 379
rect -8257 339 -8245 373
rect -6677 339 -6665 373
rect -8257 333 -6665 339
rect -6599 373 -5007 379
rect -6599 339 -6587 373
rect -5019 339 -5007 373
rect -6599 333 -5007 339
rect -4941 373 -3349 379
rect -4941 339 -4929 373
rect -3361 339 -3349 373
rect -4941 333 -3349 339
rect -3283 373 -1691 379
rect -3283 339 -3271 373
rect -1703 339 -1691 373
rect -3283 333 -1691 339
rect -1625 373 -33 379
rect -1625 339 -1613 373
rect -45 339 -33 373
rect -1625 333 -33 339
rect 33 373 1625 379
rect 33 339 45 373
rect 1613 339 1625 373
rect 33 333 1625 339
rect 1691 373 3283 379
rect 1691 339 1703 373
rect 3271 339 3283 373
rect 1691 333 3283 339
rect 3349 373 4941 379
rect 3349 339 3361 373
rect 4929 339 4941 373
rect 3349 333 4941 339
rect 5007 373 6599 379
rect 5007 339 5019 373
rect 6587 339 6599 373
rect 5007 333 6599 339
rect 6665 373 8257 379
rect 6665 339 6677 373
rect 8245 339 8257 373
rect 6665 333 8257 339
rect -8257 265 -6665 271
rect -8257 231 -8245 265
rect -6677 231 -6665 265
rect -8257 225 -6665 231
rect -6599 265 -5007 271
rect -6599 231 -6587 265
rect -5019 231 -5007 265
rect -6599 225 -5007 231
rect -4941 265 -3349 271
rect -4941 231 -4929 265
rect -3361 231 -3349 265
rect -4941 225 -3349 231
rect -3283 265 -1691 271
rect -3283 231 -3271 265
rect -1703 231 -1691 265
rect -3283 225 -1691 231
rect -1625 265 -33 271
rect -1625 231 -1613 265
rect -45 231 -33 265
rect -1625 225 -33 231
rect 33 265 1625 271
rect 33 231 45 265
rect 1613 231 1625 265
rect 33 225 1625 231
rect 1691 265 3283 271
rect 1691 231 1703 265
rect 3271 231 3283 265
rect 1691 225 3283 231
rect 3349 265 4941 271
rect 3349 231 3361 265
rect 4929 231 4941 265
rect 3349 225 4941 231
rect 5007 265 6599 271
rect 5007 231 5019 265
rect 6587 231 6599 265
rect 5007 225 6599 231
rect 6665 265 8257 271
rect 6665 231 6677 265
rect 8245 231 8257 265
rect 6665 225 8257 231
rect -8313 181 -8267 193
rect -8313 121 -8307 181
rect -8273 121 -8267 181
rect -8313 109 -8267 121
rect -6655 181 -6609 193
rect -6655 121 -6649 181
rect -6615 121 -6609 181
rect -6655 109 -6609 121
rect -4997 181 -4951 193
rect -4997 121 -4991 181
rect -4957 121 -4951 181
rect -4997 109 -4951 121
rect -3339 181 -3293 193
rect -3339 121 -3333 181
rect -3299 121 -3293 181
rect -3339 109 -3293 121
rect -1681 181 -1635 193
rect -1681 121 -1675 181
rect -1641 121 -1635 181
rect -1681 109 -1635 121
rect -23 181 23 193
rect -23 121 -17 181
rect 17 121 23 181
rect -23 109 23 121
rect 1635 181 1681 193
rect 1635 121 1641 181
rect 1675 121 1681 181
rect 1635 109 1681 121
rect 3293 181 3339 193
rect 3293 121 3299 181
rect 3333 121 3339 181
rect 3293 109 3339 121
rect 4951 181 4997 193
rect 4951 121 4957 181
rect 4991 121 4997 181
rect 4951 109 4997 121
rect 6609 181 6655 193
rect 6609 121 6615 181
rect 6649 121 6655 181
rect 6609 109 6655 121
rect 8267 181 8313 193
rect 8267 121 8273 181
rect 8307 121 8313 181
rect 8267 109 8313 121
rect -8257 71 -6665 77
rect -8257 37 -8245 71
rect -6677 37 -6665 71
rect -8257 31 -6665 37
rect -6599 71 -5007 77
rect -6599 37 -6587 71
rect -5019 37 -5007 71
rect -6599 31 -5007 37
rect -4941 71 -3349 77
rect -4941 37 -4929 71
rect -3361 37 -3349 71
rect -4941 31 -3349 37
rect -3283 71 -1691 77
rect -3283 37 -3271 71
rect -1703 37 -1691 71
rect -3283 31 -1691 37
rect -1625 71 -33 77
rect -1625 37 -1613 71
rect -45 37 -33 71
rect -1625 31 -33 37
rect 33 71 1625 77
rect 33 37 45 71
rect 1613 37 1625 71
rect 33 31 1625 37
rect 1691 71 3283 77
rect 1691 37 1703 71
rect 3271 37 3283 71
rect 1691 31 3283 37
rect 3349 71 4941 77
rect 3349 37 3361 71
rect 4929 37 4941 71
rect 3349 31 4941 37
rect 5007 71 6599 77
rect 5007 37 5019 71
rect 6587 37 6599 71
rect 5007 31 6599 37
rect 6665 71 8257 77
rect 6665 37 6677 71
rect 8245 37 8257 71
rect 6665 31 8257 37
rect -8257 -37 -6665 -31
rect -8257 -71 -8245 -37
rect -6677 -71 -6665 -37
rect -8257 -77 -6665 -71
rect -6599 -37 -5007 -31
rect -6599 -71 -6587 -37
rect -5019 -71 -5007 -37
rect -6599 -77 -5007 -71
rect -4941 -37 -3349 -31
rect -4941 -71 -4929 -37
rect -3361 -71 -3349 -37
rect -4941 -77 -3349 -71
rect -3283 -37 -1691 -31
rect -3283 -71 -3271 -37
rect -1703 -71 -1691 -37
rect -3283 -77 -1691 -71
rect -1625 -37 -33 -31
rect -1625 -71 -1613 -37
rect -45 -71 -33 -37
rect -1625 -77 -33 -71
rect 33 -37 1625 -31
rect 33 -71 45 -37
rect 1613 -71 1625 -37
rect 33 -77 1625 -71
rect 1691 -37 3283 -31
rect 1691 -71 1703 -37
rect 3271 -71 3283 -37
rect 1691 -77 3283 -71
rect 3349 -37 4941 -31
rect 3349 -71 3361 -37
rect 4929 -71 4941 -37
rect 3349 -77 4941 -71
rect 5007 -37 6599 -31
rect 5007 -71 5019 -37
rect 6587 -71 6599 -37
rect 5007 -77 6599 -71
rect 6665 -37 8257 -31
rect 6665 -71 6677 -37
rect 8245 -71 8257 -37
rect 6665 -77 8257 -71
rect -8313 -121 -8267 -109
rect -8313 -181 -8307 -121
rect -8273 -181 -8267 -121
rect -8313 -193 -8267 -181
rect -6655 -121 -6609 -109
rect -6655 -181 -6649 -121
rect -6615 -181 -6609 -121
rect -6655 -193 -6609 -181
rect -4997 -121 -4951 -109
rect -4997 -181 -4991 -121
rect -4957 -181 -4951 -121
rect -4997 -193 -4951 -181
rect -3339 -121 -3293 -109
rect -3339 -181 -3333 -121
rect -3299 -181 -3293 -121
rect -3339 -193 -3293 -181
rect -1681 -121 -1635 -109
rect -1681 -181 -1675 -121
rect -1641 -181 -1635 -121
rect -1681 -193 -1635 -181
rect -23 -121 23 -109
rect -23 -181 -17 -121
rect 17 -181 23 -121
rect -23 -193 23 -181
rect 1635 -121 1681 -109
rect 1635 -181 1641 -121
rect 1675 -181 1681 -121
rect 1635 -193 1681 -181
rect 3293 -121 3339 -109
rect 3293 -181 3299 -121
rect 3333 -181 3339 -121
rect 3293 -193 3339 -181
rect 4951 -121 4997 -109
rect 4951 -181 4957 -121
rect 4991 -181 4997 -121
rect 4951 -193 4997 -181
rect 6609 -121 6655 -109
rect 6609 -181 6615 -121
rect 6649 -181 6655 -121
rect 6609 -193 6655 -181
rect 8267 -121 8313 -109
rect 8267 -181 8273 -121
rect 8307 -181 8313 -121
rect 8267 -193 8313 -181
rect -8257 -231 -6665 -225
rect -8257 -265 -8245 -231
rect -6677 -265 -6665 -231
rect -8257 -271 -6665 -265
rect -6599 -231 -5007 -225
rect -6599 -265 -6587 -231
rect -5019 -265 -5007 -231
rect -6599 -271 -5007 -265
rect -4941 -231 -3349 -225
rect -4941 -265 -4929 -231
rect -3361 -265 -3349 -231
rect -4941 -271 -3349 -265
rect -3283 -231 -1691 -225
rect -3283 -265 -3271 -231
rect -1703 -265 -1691 -231
rect -3283 -271 -1691 -265
rect -1625 -231 -33 -225
rect -1625 -265 -1613 -231
rect -45 -265 -33 -231
rect -1625 -271 -33 -265
rect 33 -231 1625 -225
rect 33 -265 45 -231
rect 1613 -265 1625 -231
rect 33 -271 1625 -265
rect 1691 -231 3283 -225
rect 1691 -265 1703 -231
rect 3271 -265 3283 -231
rect 1691 -271 3283 -265
rect 3349 -231 4941 -225
rect 3349 -265 3361 -231
rect 4929 -265 4941 -231
rect 3349 -271 4941 -265
rect 5007 -231 6599 -225
rect 5007 -265 5019 -231
rect 6587 -265 6599 -231
rect 5007 -271 6599 -265
rect 6665 -231 8257 -225
rect 6665 -265 6677 -231
rect 8245 -265 8257 -231
rect 6665 -271 8257 -265
rect -8257 -339 -6665 -333
rect -8257 -373 -8245 -339
rect -6677 -373 -6665 -339
rect -8257 -379 -6665 -373
rect -6599 -339 -5007 -333
rect -6599 -373 -6587 -339
rect -5019 -373 -5007 -339
rect -6599 -379 -5007 -373
rect -4941 -339 -3349 -333
rect -4941 -373 -4929 -339
rect -3361 -373 -3349 -339
rect -4941 -379 -3349 -373
rect -3283 -339 -1691 -333
rect -3283 -373 -3271 -339
rect -1703 -373 -1691 -339
rect -3283 -379 -1691 -373
rect -1625 -339 -33 -333
rect -1625 -373 -1613 -339
rect -45 -373 -33 -339
rect -1625 -379 -33 -373
rect 33 -339 1625 -333
rect 33 -373 45 -339
rect 1613 -373 1625 -339
rect 33 -379 1625 -373
rect 1691 -339 3283 -333
rect 1691 -373 1703 -339
rect 3271 -373 3283 -339
rect 1691 -379 3283 -373
rect 3349 -339 4941 -333
rect 3349 -373 3361 -339
rect 4929 -373 4941 -339
rect 3349 -379 4941 -373
rect 5007 -339 6599 -333
rect 5007 -373 5019 -339
rect 6587 -373 6599 -339
rect 5007 -379 6599 -373
rect 6665 -339 8257 -333
rect 6665 -373 6677 -339
rect 8245 -373 8257 -339
rect 6665 -379 8257 -373
rect -8313 -423 -8267 -411
rect -8313 -483 -8307 -423
rect -8273 -483 -8267 -423
rect -8313 -495 -8267 -483
rect -6655 -423 -6609 -411
rect -6655 -483 -6649 -423
rect -6615 -483 -6609 -423
rect -6655 -495 -6609 -483
rect -4997 -423 -4951 -411
rect -4997 -483 -4991 -423
rect -4957 -483 -4951 -423
rect -4997 -495 -4951 -483
rect -3339 -423 -3293 -411
rect -3339 -483 -3333 -423
rect -3299 -483 -3293 -423
rect -3339 -495 -3293 -483
rect -1681 -423 -1635 -411
rect -1681 -483 -1675 -423
rect -1641 -483 -1635 -423
rect -1681 -495 -1635 -483
rect -23 -423 23 -411
rect -23 -483 -17 -423
rect 17 -483 23 -423
rect -23 -495 23 -483
rect 1635 -423 1681 -411
rect 1635 -483 1641 -423
rect 1675 -483 1681 -423
rect 1635 -495 1681 -483
rect 3293 -423 3339 -411
rect 3293 -483 3299 -423
rect 3333 -483 3339 -423
rect 3293 -495 3339 -483
rect 4951 -423 4997 -411
rect 4951 -483 4957 -423
rect 4991 -483 4997 -423
rect 4951 -495 4997 -483
rect 6609 -423 6655 -411
rect 6609 -483 6615 -423
rect 6649 -483 6655 -423
rect 6609 -495 6655 -483
rect 8267 -423 8313 -411
rect 8267 -483 8273 -423
rect 8307 -483 8313 -423
rect 8267 -495 8313 -483
rect -8257 -533 -6665 -527
rect -8257 -567 -8245 -533
rect -6677 -567 -6665 -533
rect -8257 -573 -6665 -567
rect -6599 -533 -5007 -527
rect -6599 -567 -6587 -533
rect -5019 -567 -5007 -533
rect -6599 -573 -5007 -567
rect -4941 -533 -3349 -527
rect -4941 -567 -4929 -533
rect -3361 -567 -3349 -533
rect -4941 -573 -3349 -567
rect -3283 -533 -1691 -527
rect -3283 -567 -3271 -533
rect -1703 -567 -1691 -533
rect -3283 -573 -1691 -567
rect -1625 -533 -33 -527
rect -1625 -567 -1613 -533
rect -45 -567 -33 -533
rect -1625 -573 -33 -567
rect 33 -533 1625 -527
rect 33 -567 45 -533
rect 1613 -567 1625 -533
rect 33 -573 1625 -567
rect 1691 -533 3283 -527
rect 1691 -567 1703 -533
rect 3271 -567 3283 -533
rect 1691 -573 3283 -567
rect 3349 -533 4941 -527
rect 3349 -567 3361 -533
rect 4929 -567 4941 -533
rect 3349 -573 4941 -567
rect 5007 -533 6599 -527
rect 5007 -567 5019 -533
rect 6587 -567 6599 -533
rect 5007 -573 6599 -567
rect 6665 -533 8257 -527
rect 6665 -567 6677 -533
rect 8245 -567 8257 -533
rect 6665 -573 8257 -567
<< properties >>
string FIXED_BBOX -8424 -688 8424 688
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 8.0 m 4 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
