* NGSPICE file created from overvoltage_ana_rcx.ext - technology: sky130A

.subckt overvoltage_ana_rcx otrip_decoded[14] otrip_decoded[13] otrip_decoded[11]
+ otrip_decoded[10] otrip_decoded[1] otrip_decoded[0] ena itest ibg_200n otrip_decoded[7]
+ otrip_decoded[4] vbg_1v2 vin isrc_sel otrip_decoded[5] otrip_decoded[8] otrip_decoded[2]
+ ovout otrip_decoded[15] otrip_decoded[9] otrip_decoded[12] otrip_decoded[3] otrip_decoded[6]
+ avss dvdd dvss avdd
X0 rstring_mux_0.vtrip12.t4 rstring_mux_0.otrip_decoded_avdd[12] vin.t27 avss.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 comparator_0.vt comparator_0.vn avss.t193 avss.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2 comparator_0.vt vin.t94 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X3 rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y rstring_mux_0.otrip_decoded_avdd[15] avss.t151 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X4 a_5346_n3990# a_4921_n3946# dvss.t223 dvss.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X5 avdd.t196 a_429_n2876# a_1122_n3990# avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X6 avss.t146 avss.t145 avss.t146 avss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X7 dvss.t206 otrip_decoded[0].t0 a_n8119_n2964# dvss.t205 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X8 a_n18769_n11914# a_n18391_n15834# avss.t147 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X9 avdd.t35 comparator_0.vpp comparator_0.vpp avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X10 rstring_mux_0.vtrip9.t2 rstring_mux_0.vtrip8.t2 avss.t246 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X11 vin.t42 avdd.t179 vin.t42 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X12 rstring_mux_0.otrip_decoded_b_avdd[1] rstring_mux_0.otrip_decoded_avdd[1] avss.t374 avss.t373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X13 dvss.t134 a_7033_n3946# a_7458_n3990# dvss.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X14 avdd.t34 comparator_0.vpp comparator_0.vnn avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X15 rstring_mux_0.otrip_decoded_avdd[5] a_n2588_n1478# avdd.t215 avdd.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X16 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t4 dvdd.t73 dvdd.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_7458_n3990# a_7033_n3946# dvss.t132 dvss.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X18 ibias_gen_0.vr.t1 ibias_gen_0.vn0.t19 ibias_gen_0.vp0.t1 avss.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X19 avdd.t291 a_2541_n2876# a_3234_n3990# avdd.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X20 a_n26830_n2937# a_n27208_n10337# avss.t309 sky130_fd_pr__res_xhigh_po_1p41 l=35
X21 comparator_0.vt vin.t95 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X22 dvss.t45 a_9145_n3946# a_9570_n3990# dvss.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X23 dvss.t178 sky130_fd_sc_hd__inv_4_0.Y ovout.t15 dvss.t177 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 rstring_mux_0.otrip_decoded_avdd[8] a_1636_n3212# dvss.t124 dvss.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X25 dvss.t237 a_6765_n2876# a_7972_n3212# dvss.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X26 avdd.t205 ibias_gen_0.isrc_sel ibias_gen_0.isrc_sel_b avdd.t204 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X27 a_n8951_9395# a_n8573_1995# avss.t361 sky130_fd_pr__res_xhigh_po_1p41 l=35
X28 dvdd.t59 sky130_fd_sc_hd__inv_4_0.Y ovout.t31 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 itest.t1 ibias_gen_0.vp.t7 avdd.t45 avdd.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X30 vin.t41 avdd.t177 vin.t41 avdd.t178 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X31 a_n24562_n2937# a_n24184_n10337# avss.t177 sky130_fd_pr__res_xhigh_po_1p41 l=35
X32 a_n21538_n2937# a_n21160_n10337# avss.t339 sky130_fd_pr__res_xhigh_po_1p41 l=35
X33 avdd.t259 a_4653_n2876# a_5346_n3990# avdd.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X34 vin.t40 avdd.t175 vin.t40 avdd.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X35 rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.otrip_decoded_avdd[2] avss.t241 avss.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X36 avss.t327 ibias_gen_0.ena rstring_mux_0.ena_b avss.t326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X37 avdd.t174 avdd.t173 avdd.t174 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=8
X38 a_n26830_n2937# a_n26452_n10337# avss.t59 sky130_fd_pr__res_xhigh_po_1p41 l=35
X39 a_n23806_n2937# a_n23428_n10337# avss.t307 sky130_fd_pr__res_xhigh_po_1p41 l=35
X40 rstring_mux_0.vtrip10.t1 rstring_mux_0.otrip_decoded_avdd[10] vin.t3 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X41 dcomp comparator_0.n1 avss.t41 avss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X42 a_n7326_n3990# a_n7751_n3946# dvss.t486 dvss.t485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X43 rstring_mux_0.otrip_decoded_avdd[10] a_3748_n3212# dvss.t271 dvss.t270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X44 comparator_0.vpp vin.t96 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X45 schmitt_trigger_0.out.t0 schmitt_trigger_0.m.t14 dvdd.t103 dvdd.t102 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X46 avdd.t353 a_n3795_n1142# a_n2588_n1478# avdd.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X47 a_9203_n11914# a_9581_n15834# avss.t376 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X48 ibias_gen_0.vp1.t16 ibias_gen_0.vp1.t15 avdd.t424 avdd.t423 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X49 a_n15529_n2223# ibias_gen_0.isrc_sel_b ibias_gen_0.vn1.t9 avdd.t428 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X50 a_n1683_n1142# a_n1783_n1230# dvss.t541 dvss.t540 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X51 dvss.t319 otrip_decoded[11].t0 a_2441_n1230# dvss.t318 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X52 avdd.t11 a_n3102_n2256# a_n3795_n1142# avdd.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X53 a_2809_n3946# a_2441_n2964# dvdd.t91 dvdd.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X54 avdd.t252 a_6765_n2876# a_7458_n3990# avdd.t251 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X55 dcomp comparator_0.n1 avdd.t67 avdd.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X56 comparator_0.vt vbg_1v2.t0 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X57 a_n6673_n11914# a_n6295_n15834# avss.t331 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X58 rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.otrip_decoded_avdd[6] avdd.t217 avdd.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X59 rstring_mux_0.vtrip11.t3 rstring_mux_0.otrip_decoded_b_avdd[11] vin.t51 avdd.t312 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X60 ibias_gen_0.vn0.t7 vbg_1v2.t1 ibias_gen_0.vstart.t10 avss.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X61 ibias_gen_0.vr.t4 a_n20404_n10337# avss.t218 sky130_fd_pr__res_xhigh_po_1p41 l=35
X62 avdd.t327 a_n5907_n1142# a_n4700_n1478# avdd.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X63 comparator_0.vpp comparator_0.vnn avdd.t237 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X64 a_n13487_9395# a_n13109_1995# avss.t251 sky130_fd_pr__res_xhigh_po_1p41 l=35
X65 dvdd.t71 schmitt_trigger_0.out.t5 sky130_fd_sc_hd__inv_4_0.Y dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X66 a_n3795_n1142# a_n3895_n1230# dvss.t146 dvss.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X67 a_2541_n1142# a_2441_n1230# dvss.t269 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X68 a_7033_n3946# a_6665_n2964# dvdd.t119 dvdd.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X69 avdd.t236 comparator_0.vnn comparator_0.vpp avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X70 avdd.t172 avdd.t170 avdd.t171 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=8
X71 avdd.t169 avdd.t168 avdd.t169 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=8
X72 ovout.t30 sky130_fd_sc_hd__inv_4_0.Y dvdd.t57 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X73 rstring_mux_0.vtrip5.t4 rstring_mux_0.vtrip4.t3 avss.t340 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X74 a_n14243_9395# a_n14621_1995# avss.t207 sky130_fd_pr__res_xhigh_po_1p41 l=35
X75 dvdd.t101 otrip_decoded[6].t0 a_n1783_n2964# dvdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X76 dvss.t435 a_8877_n1142# a_10084_n1478# dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X77 rstring_mux_0.otrip_decoded_avdd[13] a_5860_n1478# avdd.t188 avdd.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X78 a_n25573_n11914# a_n25195_n15834# avss.t47 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X79 rstring_mux_0.otrip_decoded_b_avdd[1] rstring_mux_0.otrip_decoded_avdd[1] avdd.t438 avdd.t437 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X80 dvss.t307 a_2541_n2876# a_3748_n3212# dvss.t306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X81 comparator_0.vm comparator_0.vm avss.t250 avss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X82 comparator_0.vnn comparator_0.vpp avdd.t33 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X83 avdd.t235 comparator_0.vnn comparator_0.vnn avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X84 comparator_0.vt vbg_1v2.t2 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X85 avdd.t383 a_n8019_n1142# a_n6812_n1478# avdd.t206 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X86 a_n9697_n11914# a_n10075_n15834# avss.t357 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X87 vin.t7 rstring_mux_0.otrip_decoded_b_avdd[13] rstring_mux_0.vtrip13.t1 avdd.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X88 rstring_mux_0.otrip_decoded_avdd[5] a_n2588_n1478# dvss.t180 dvss.t179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X89 schmitt_trigger_0.m.t0 schmitt_trigger_0.in.t1 dvdd.t15 dvdd.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X90 a_4653_n1142# a_4553_n1230# dvss.t521 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X91 a_9145_n3946# a_8777_n2964# dvdd.t89 dvdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X92 a_n13477_n11914# a_n13099_n15834# avss.t198 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X93 dvdd.t139 otrip_decoded[4].t0 a_n3895_n2964# dvdd.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X94 a_n11975_9395# a_n11597_1995# avss.t345 sky130_fd_pr__res_xhigh_po_1p41 l=35
X95 dvss.t514 otrip_decoded[9].t0 a_329_n1230# dvss.t513 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X96 a_697_n3946# a_329_n2964# dvdd.t75 dvdd.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X97 comparator_0.n1 comparator_0.n0 avdd.t247 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X98 a_n20281_n11914# a_n20659_n15834# avss.t380 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X99 avdd.t65 comparator_0.n1 dcomp avdd.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X100 avdd.t275 a_429_n1142# a_1636_n1478# avdd.t274 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X101 avdd.t416 rstring_mux_0.ena_b rstring_mux_0.vtop.t16 avdd.t415 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X102 dvss.t249 a_4653_n2876# a_5860_n3212# dvss.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X103 a_n5161_n11914# a_n4783_n15834# avss.t298 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X104 comparator_0.n1 comparator_0.n0 avss.t212 avss.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X105 comparator_0.vpp vin.t97 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X106 ovout.t29 sky130_fd_sc_hd__inv_4_0.Y dvdd.t55 dvdd.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X107 dvss.t176 sky130_fd_sc_hd__inv_4_0.Y ovout.t14 dvss.t175 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X108 ibias_gen_0.vp0.t5 ibias_gen_0.vp0.t4 avdd.t365 avdd.t364 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X109 rstring_mux_0.otrip_decoded_avdd[3] a_n4700_n1478# dvss.t63 dvss.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X110 schmitt_trigger_0.m.t1 schmitt_trigger_0.in.t2 dvss.t112 dvss.t111 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X111 a_6765_n1142# a_6665_n1230# dvss.t92 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X112 a_n5161_n11914# a_n5539_n15834# avss.t19 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X113 dvss.t430 dvss.t428 schmitt_trigger_0.m.t12 dvss.t429 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X114 rstring_mux_0.vtop.t15 rstring_mux_0.ena_b avdd.t414 avdd.t413 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X115 ibias_gen_0.ena_b ibias_gen_0.ena avss.t325 avss.t324 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X116 rstring_mux_0.otrip_decoded_avdd[2] a_n4700_n3212# avdd.t418 avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X117 vin.t86 rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.vtrip6.t5 avdd.t436 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X118 dvdd.t126 otrip_decoded[2].t0 a_n6007_n2964# dvdd.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X119 avss.t144 avss.t142 avss.t143 avss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X120 dcomp comparator_0.n1 avdd.t63 avdd.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X121 comparator_0.vnn comparator_0.vpp avdd.t32 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X122 avdd.t31 comparator_0.vpp comparator_0.n0 avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X123 ibias_gen_0.vp.t4 ibias_gen_0.ena avdd.t347 avdd.t346 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X124 avdd.t283 a_1122_n2256# a_429_n1142# avdd.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X125 avdd.t412 rstring_mux_0.ena_b rstring_mux_0.vtop.t14 avdd.t411 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X126 avdd.t47 ibias_gen_0.vp.t8 ibias_gen_0.ibias avdd.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X127 rstring_mux_0.otrip_decoded_b_avdd[8] rstring_mux_0.otrip_decoded_avdd[8] avss.t158 avss.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X128 comparator_0.vpp ibias_gen_0.ena avdd.t345 avdd.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X129 ibias_gen_0.vn0.t4 ibias_gen_0.vn0.t3 ibias_gen_0.ve.t1 avss.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X130 ibias_gen_0.vp.t5 ibias_gen_0.isrc_sel_b ibias_gen_0.vp0.t10 avss.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X131 vin.t39 avdd.t166 vin.t39 avdd.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X132 dvss.t174 sky130_fd_sc_hd__inv_4_0.Y ovout.t13 dvss.t173 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X133 rstring_mux_0.vtop.t13 rstring_mux_0.ena_b avdd.t410 avdd.t409 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X134 ibias_gen_0.vp1.t4 ibias_gen_0.vn1.t10 avss.t287 avss.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X135 a_n24061_n11914# a_n23683_n15834# avss.t301 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X136 comparator_0.vn ibias_gen_0.ena ibias_gen_0.ibias avss.t323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X137 a_n7751_n2212# a_n8119_n1230# dvss.t104 dvss.t103 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X138 rstring_mux_0.otrip_decoded_avdd[0] a_n6812_n3212# avdd.t269 avdd.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X139 rstring_mux_0.otrip_decoded_b_avdd[12] rstring_mux_0.otrip_decoded_avdd[12] avss.t234 avss.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X140 comparator_0.vnn ibias_gen_0.ena avdd.t343 avdd.t342 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X141 a_n24061_n11914# a_n24439_n15834# avss.t219 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X142 dvdd.t5 otrip_decoded[0].t1 a_n8119_n2964# dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X143 a_9959_n11914# a_10337_n15834# avss.t154 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X144 vin.t48 rstring_mux_0.otrip_decoded_b_avdd[1] rstring_mux_0.vtrip1.t1 avdd.t302 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X145 rstring_mux_0.otrip_decoded_avdd[9] a_1636_n1478# avdd.t350 avdd.t274 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X146 avdd.t380 a_6765_n1142# a_7972_n1478# avdd.t379 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X147 avdd.t254 a_3234_n2256# a_2541_n1142# avdd.t253 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X148 a_n8195_9395# schmitt_trigger_0.in.t0 avss.t274 sky130_fd_pr__res_xhigh_po_1p41 l=35
X149 a_n11965_n11914# a_n11587_n15834# avss.t185 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X150 a_n8941_n11914# a_n8563_n15834# avss.t48 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X151 a_3911_n11914# a_4289_n15834# avss.t4 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X152 vin.t70 rstring_mux_0.otrip_decoded_avdd[0] rstring_mux_0.vtrip0.t5 avss.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X153 dvss.t114 schmitt_trigger_0.in.t3 schmitt_trigger_0.m.t2 dvss.t113 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X154 a_n8951_9395# a_n9329_1995# avss.t153 sky130_fd_pr__res_xhigh_po_1p41 l=35
X155 avss.t141 avss.t139 avss.t140 avss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X156 vin.t75 avdd.t164 vin.t75 avdd.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X157 comparator_0.vpp comparator_0.vpp avdd.t30 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X158 dvdd.t87 otrip_decoded[11].t1 a_2441_n1230# dvdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X159 vin.t74 avdd.t162 vin.t74 avdd.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X160 rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.otrip_decoded_avdd[4] avss.t52 avss.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X161 avdd.t49 ibias_gen_0.vp.t9 itest.t0 avdd.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X162 vin.t9 rstring_mux_0.otrip_decoded_avdd[4] rstring_mux_0.vtrip4.t2 avss.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X163 ibias_gen_0.vstart.t9 vbg_1v2.t3 ibias_gen_0.vn0.t8 avss.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X164 comparator_0.ena_b ibias_gen_0.ena avdd.t341 avdd.t340 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X165 ibias_gen_0.isrc_sel_b avss.t137 ibias_gen_0.ena_b avss.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X166 a_n1683_n1142# a_n1783_n1230# dvss.t539 dvss.t538 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X167 a_n20782_n2937# a_n21160_n10337# avss.t206 sky130_fd_pr__res_xhigh_po_1p41 l=35
X168 avdd.t234 comparator_0.vnn comparator_0.vpp avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X169 rstring_mux_0.otrip_decoded_avdd[11] a_3748_n1478# avdd.t324 avdd.t318 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X170 avdd.t161 avdd.t160 avdd.t161 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=8
X171 dvdd.t17 schmitt_trigger_0.in.t4 schmitt_trigger_0.m.t3 dvdd.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X172 avdd.t249 a_5346_n2256# a_4653_n1142# avdd.t248 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X173 comparator_0.vn comparator_0.ena_b ibias_gen_0.ibias avdd.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X174 ovout.t28 sky130_fd_sc_hd__inv_4_0.Y dvdd.t53 dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X175 a_n27841_n11914# a_n27463_n15834# avss.t341 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X176 rstring_mux_0.vtop.t12 rstring_mux_0.ena_b avdd.t408 avdd.t407 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X177 a_n3795_n1142# a_n3895_n1230# dvss.t144 dvss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X178 a_n14989_n11914# a_n15367_n15834# avss.t346 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X179 rstring_mux_0.vtrip13.t0 rstring_mux_0.otrip_decoded_b_avdd[13] vin.t6 avdd.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X180 comparator_0.vnn avss.t385 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X181 avdd.t422 ibias_gen_0.vp1.t13 ibias_gen_0.vp1.t14 avdd.t421 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X182 dvss.t172 sky130_fd_sc_hd__inv_4_0.Y ovout.t12 dvss.t171 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X183 vin.t82 rstring_mux_0.otrip_decoded_avdd[11] rstring_mux_0.vtrip11.t5 avss.t369 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X184 a_7691_n11914# a_8069_n15834# avss.t271 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X185 rstring_mux_0.vtrip3.t1 rstring_mux_0.otrip_decoded_avdd[3] vin.t1 avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X186 vin.t92 rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y rstring_mux_0.vtrip15.t5 avdd.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X187 a_n15745_n11914# a_n15367_n15834# avss.t213 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X188 dvss.t498 a_n6007_n1230# a_n5907_n1142# dvss.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X189 dvss.t520 a_4553_n1230# a_4653_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X190 comparator_0.vpp vin.t98 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X191 avss.t288 ibias_gen_0.vn1.t11 ibias_gen_0.vp1.t5 avss.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X192 ovout.t27 sky130_fd_sc_hd__inv_4_0.Y dvdd.t51 dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X193 avdd.t304 a_7458_n2256# a_6765_n1142# avdd.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X194 rstring_mux_0.vtrip9.t1 rstring_mux_0.otrip_decoded_avdd[9] vin.t23 avss.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X195 rstring_mux_0.vtrip0.t4 rstring_mux_0.otrip_decoded_avdd[0] vin.t69 avss.t349 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X196 ibias_gen_0.vp1.t6 ibias_gen_0.vn1.t12 avss.t289 avss.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X197 rstring_mux_0.otrip_decoded_avdd[14] a_7972_n3212# avdd.t73 avdd.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X198 ibias_gen_0.vp.t2 ibias_gen_0.isrc_sel ibias_gen_0.vp0.t8 avdd.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X199 comparator_0.vt vbg_1v2.t4 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X200 a_n5907_n1142# a_n6007_n1230# dvss.t496 dvss.t495 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X201 rstring_mux_0.vtrip15.t3 a_2777_n15834# avss.t256 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X202 avdd.t29 comparator_0.vpp comparator_0.vpp avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X203 avss.t290 ibias_gen_0.vn1.t13 ibias_gen_0.vp1.t7 avss.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X204 rstring_mux_0.vtrip4.t1 rstring_mux_0.otrip_decoded_avdd[4] vin.t8 avss.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X205 avdd.t159 avdd.t158 avdd.t159 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X206 dvss.t170 sky130_fd_sc_hd__inv_4_0.Y ovout.t11 dvss.t169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X207 dvdd.t1 otrip_decoded[9].t1 a_329_n1230# dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X208 vin.t29 rstring_mux_0.otrip_decoded_avdd[2] rstring_mux_0.vtrip2.t1 avss.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X209 a_n14999_9395# a_n14621_1995# avss.t220 sky130_fd_pr__res_xhigh_po_1p41 l=35
X210 a_3155_n11914# a_2777_n15834# avss.t344 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X211 vin.t52 rstring_mux_0.otrip_decoded_b_avdd[11] rstring_mux_0.vtrip11.t2 avdd.t311 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X212 avdd.t319 a_2541_n1142# a_3748_n1478# avdd.t318 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X213 a_n10453_n11914# a_n10831_n15834# avss.t23 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X214 rstring_mux_0.vtrip8.t1 rstring_mux_0.otrip_decoded_avdd[8] vin.t12 avss.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X215 rstring_mux_0.vtrip7.t2 rstring_mux_0.otrip_decoded_avdd[7] vin.t37 avss.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X216 a_n10463_9395# a_n10085_1995# avss.t21 sky130_fd_pr__res_xhigh_po_1p41 l=35
X217 dvss.t102 a_n8119_n1230# a_n8019_n1142# dvss.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X218 dvss.t91 a_6665_n1230# a_6765_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X219 avdd.t261 a_9570_n2256# a_8877_n1142# avdd.t260 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X220 vin.t73 avdd.t156 vin.t73 avdd.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X221 vin.t46 avss.t135 vin.t46 avss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X222 comparator_0.vnn comparator_0.vnn avdd.t233 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X223 avdd.t155 avdd.t153 avdd.t155 avdd.t154 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X224 dvss.t281 a_697_n2212# a_1122_n2256# dvss.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X225 a_8877_n1142# a_8777_n1230# dvss.t83 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X226 a_n18769_n11914# a_n19147_n15834# avss.t236 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X227 ibias_gen_0.vp.t1 avss.t133 ibias_gen_0.vp.t1 avss.t134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X228 rstring_mux_0.vtrip9.t5 rstring_mux_0.vtrip10.t5 avss.t384 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X229 avss.t191 comparator_0.vn comparator_0.vn avss.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X230 comparator_0.vpp vin.t99 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X231 a_n19525_n11914# a_n19147_n15834# avss.t208 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X232 dvss.t194 a_8877_n2876# a_10084_n3212# dvss.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X233 a_429_n1142# a_329_n1230# dvss.t213 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X234 rstring_mux_0.otrip_decoded_avdd[6] a_n476_n3212# avdd.t71 avdd.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X235 a_n26329_n11914# a_n25951_n15834# avss.t245 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X236 a_n11975_9395# a_n12353_1995# avss.t46 sky130_fd_pr__res_xhigh_po_1p41 l=35
X237 avdd.t288 a_4653_n1142# a_5860_n1478# avdd.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X238 comparator_0.vpp comparator_0.vnn avdd.t232 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X239 dvss.t82 a_8777_n1230# a_8877_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X240 vin.t80 rstring_mux_0.otrip_decoded_avdd[13] rstring_mux_0.vtrip13.t5 avss.t365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X241 avdd.t427 ibias_gen_0.isrc_sel_b ibias_gen_0.vp0.t11 avdd.t426 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X242 vin.t72 avdd.t151 vin.t72 avdd.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X243 rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.otrip_decoded_avdd[0] avss.t348 avss.t347 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X244 comparator_0.vm comparator_0.ena_b avss.t184 avss.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X245 rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.otrip_decoded_avdd[4] avdd.t69 avdd.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X246 ovout.t26 sky130_fd_sc_hd__inv_4_0.Y dvdd.t49 dvdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X247 a_6179_n11914# a_6557_n15834# avss.t270 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X248 dcomp comparator_0.n1 avss.t39 avss.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X249 dvss.t212 a_329_n1230# a_429_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X250 a_n14233_n11914# a_n13855_n15834# avss.t57 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X251 rstring_mux_0.vtrip5.t1 rstring_mux_0.otrip_decoded_avdd[5] vin.t19 avss.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X252 avdd.t363 ibias_gen_0.vp0.t2 ibias_gen_0.vp0.t3 avdd.t362 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X253 a_8877_n1142# a_8777_n1230# dvss.t81 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X254 a_n7751_n2212# a_n8119_n1230# dvdd.t11 dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X255 vin.t56 rstring_mux_0.otrip_decoded_b_avdd[10] rstring_mux_0.vtrip10.t4 avdd.t323 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X256 a_n14233_n11914# a_n14611_n15834# avss.t231 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X257 ibias_gen_0.vn0.t9 vbg_1v2.t5 ibias_gen_0.vstart.t8 avss.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X258 a_5346_n2256# a_4921_n2212# dvss.t470 dvss.t469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X259 avdd.t231 comparator_0.vnn comparator_0.vnn avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X260 comparator_0.n0 comparator_0.vpp avdd.t28 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X261 avdd.t202 ibias_gen_0.isrc_sel a_n16775_n2223# avdd.t201 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X262 schmitt_trigger_0.m.t11 schmitt_trigger_0.out.t6 dvdd.t69 dvdd.t68 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X263 rstring_mux_0.vtrip2.t0 rstring_mux_0.otrip_decoded_avdd[2] vin.t28 avss.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X264 dvdd.t105 schmitt_trigger_0.m.t15 schmitt_trigger_0.out.t1 dvdd.t104 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X265 comparator_0.vpp vin.t100 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X266 rstring_mux_0.vtrip13.t3 rstring_mux_0.vtrip12.t5 avss.t264 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X267 avdd.t339 ibias_gen_0.ena ibias_gen_0.vp1.t12 avdd.t338 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X268 ovout.t25 sky130_fd_sc_hd__inv_4_0.Y dvdd.t47 dvdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X269 ibias_gen_0.vp1.t2 ibias_gen_0.isrc_sel avdd.t200 avdd.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X270 rstring_mux_0.vtrip6.t4 rstring_mux_0.otrip_decoded_b_avdd[6] vin.t85 avdd.t435 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X271 ibias_gen_0.ena a_10084_n3212# dvss.t460 dvss.t459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X272 rstring_mux_0.vtrip13.t2 rstring_mux_0.vtrip14.t0 avss.t53 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X273 comparator_0.vt vbg_1v2.t6 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X274 a_7458_n2256# a_7033_n2212# dvss.t247 dvss.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X275 avdd.t76 a_n1683_n2876# a_n476_n3212# avdd.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X276 vin.t45 avss.t131 vin.t45 avss.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X277 a_9959_n11914# a_9581_n15834# avss.t337 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X278 avdd.t295 a_n990_n3990# a_n1683_n2876# avdd.t294 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X279 a_n1683_n2876# a_n1783_n2964# dvss.t399 dvss.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X280 dvss.t363 otrip_decoded[10].t0 a_2441_n2964# dvss.t362 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X281 a_n18013_n11914# a_n17635_n15834# avss.t225 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X282 vin.t44 avss.t129 vin.t44 avss.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X283 a_2541_n1142# a_2441_n1230# dvss.t268 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X284 a_n990_n2256# a_n1415_n2212# dvss.t13 dvss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X285 a_n18013_n11914# a_n18391_n15834# avss.t176 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X286 a_n3795_n1142# a_n3895_n1230# dvss.t142 dvss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X287 dvss.t450 a_n1683_n1142# a_n476_n1478# dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X288 avdd.t190 a_n5214_n2256# a_n5907_n1142# avdd.t189 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X289 vin.t43 avss.t127 vin.t43 avss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X290 rstring_mux_0.vtrip1.t0 rstring_mux_0.otrip_decoded_b_avdd[1] vin.t47 avdd.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X291 ibias_gen_0.vp.t0 avdd.t149 ibias_gen_0.vp.t0 avdd.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X292 comparator_0.vnn avss.t386 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X293 dvss.t168 sky130_fd_sc_hd__inv_4_0.Y ovout.t10 dvss.t167 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X294 dvss.t457 a_n8019_n1142# a_n6812_n1478# dvss.t456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X295 dvss.t267 a_2441_n1230# a_2541_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X296 rstring_mux_0.otrip_decoded_b_avdd[5] rstring_mux_0.otrip_decoded_avdd[5] avss.t202 avss.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X297 a_n3795_n2876# a_n3895_n2964# dvss.t235 dvss.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X298 a_2541_n2876# a_2441_n2964# dvss.t343 dvss.t342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X299 a_n12721_n11914# a_n13099_n15834# avss.t379 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X300 a_5423_n11914# a_5045_n15834# avss.t257 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X301 a_n26074_n2937# a_n26452_n10337# avss.t15 sky130_fd_pr__res_xhigh_po_1p41 l=35
X302 a_n23050_n2937# a_n23428_n10337# avss.t329 sky130_fd_pr__res_xhigh_po_1p41 l=35
X303 dvss.t262 a_10515_n2156# a_10874_n2222# dvss.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X304 rstring_mux_0.vtrip3.t2 rstring_mux_0.vtrip4.t0 avss.t16 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X305 a_n5907_n1142# a_n6007_n1230# dvss.t494 dvss.t493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X306 rstring_mux_0.otrip_decoded_avdd[11] a_3748_n1478# dvss.t385 dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X307 a_n5907_n1142# a_n6007_n1230# dvss.t492 dvss.t491 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X308 a_4653_n1142# a_4553_n1230# dvss.t519 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X309 avdd.t329 a_n7326_n2256# a_n8019_n1142# avdd.t328 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X310 rstring_mux_0.vtrip3.t5 rstring_mux_0.vtrip2.t4 avss.t375 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X311 avdd.t148 avdd.t146 avdd.t147 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=8
X312 a_n25318_n2937# a_n25696_n10337# avss.t305 sky130_fd_pr__res_xhigh_po_1p41 l=35
X313 ibias_gen_0.vn1.t7 ibias_gen_0.vn1.t6 avss.t286 avss.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X314 dvss.t317 a_10515_n1026# a_10515_n2156# dvss.t316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X315 a_n1415_n2212# a_n1783_n1230# dvss.t537 dvss.t536 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X316 dvss.t100 a_n8119_n1230# a_n8019_n1142# dvss.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X317 dvdd.t67 schmitt_trigger_0.out.t7 sky130_fd_sc_hd__inv_4_0.Y dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X318 a_4653_n2876# a_4553_n2964# dvss.t411 dvss.t410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X319 comparator_0.vpp comparator_0.vnn avdd.t230 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X320 avss.t126 avss.t124 avss.t125 avss.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X321 schmitt_trigger_0.m.t8 schmitt_trigger_0.out.t8 dvss.t345 dvss.t344 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X322 avdd.t229 comparator_0.vnn comparator_0.vpp avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X323 comparator_0.vnn avss.t387 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X324 a_n8019_n1142# a_n8119_n1230# dvss.t98 dvss.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X325 a_6765_n1142# a_6665_n1230# dvss.t90 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X326 dvss.t437 isrc_sel.t0 a_8777_n1230# dvss.t436 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X327 a_n21037_n11914# a_n20659_n15834# avss.t314 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X328 rstring_mux_0.vtrip2.t3 rstring_mux_0.otrip_decoded_b_avdd[2] vin.t62 avdd.t376 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X329 avdd.t145 avdd.t144 avdd.t145 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=8
X330 a_n14999_9395# vl.t0 avss.t6 sky130_fd_pr__res_xhigh_po_1p41 l=35
X331 a_n8019_n1142# a_n8119_n1230# dvss.t96 dvss.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X332 rstring_mux_0.otrip_decoded_b_avdd[7] rstring_mux_0.otrip_decoded_avdd[7] avss.t268 avss.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X333 rstring_mux_0.otrip_decoded_b_avdd[14] rstring_mux_0.otrip_decoded_avdd[14] avdd.t267 avdd.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X334 dvss.t25 otrip_decoded[8].t0 a_329_n2964# dvss.t24 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X335 a_n3527_n2212# a_n3895_n1230# dvss.t140 dvss.t139 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X336 rstring_mux_0.otrip_decoded_avdd[4] a_n2588_n3212# avdd.t443 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X337 a_n21037_n11914# a_n21415_n15834# avss.t308 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X338 a_8447_n11914# a_8825_n15834# avss.t237 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X339 ovout.t24 sky130_fd_sc_hd__inv_4_0.Y dvdd.t45 dvdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X340 a_429_n1142# a_329_n1230# dvss.t211 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X341 vin.t36 avss.t122 vin.t36 avss.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X342 rstring_mux_0.vtrip10.t3 rstring_mux_0.otrip_decoded_b_avdd[10] vin.t55 avdd.t322 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X343 avss.t37 comparator_0.n1 dcomp avss.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X344 a_n16501_n11914# a_n16879_n15834# avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X345 a_9203_n11914# a_8825_n15834# avss.t306 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X346 a_n10463_9395# a_n10841_1995# avss.t42 sky130_fd_pr__res_xhigh_po_1p41 l=35
X347 ibias_gen_0.vp1.t8 ibias_gen_0.vn1.t14 avss.t291 avss.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X348 a_n5917_n11914# a_n5539_n15834# avss.t56 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X349 rstring_mux_0.otrip_decoded_b_avdd[14] rstring_mux_0.otrip_decoded_avdd[14] avss.t229 avss.t228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X350 a_6765_n2876# a_6665_n2964# dvss.t427 dvss.t426 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X351 ibias_gen_0.vp0.t6 avdd.t141 avdd.t143 avdd.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X352 dvss.t375 a_2809_n2212# a_3234_n2256# dvss.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X353 comparator_0.vt vbg_1v2.t7 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X354 dvss.t210 a_329_n1230# a_429_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X355 dvdd.t133 a_10874_n2222# vl.t2 dvdd.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X356 avss.t121 avss.t119 ibias_gen_0.vr.t3 avss.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X357 avdd.t361 a_8877_n1142# a_10084_n1478# avdd.t360 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X358 avdd.t61 comparator_0.n1 dcomp avdd.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X359 a_3911_n11914# a_3533_n15834# avss.t333 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X360 a_n5639_n2212# a_n6007_n1230# dvss.t490 dvss.t489 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X361 vin.t71 avdd.t139 vin.t71 avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X362 dcomp comparator_0.n1 avss.t35 avss.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X363 comparator_0.vnn vbg_1v2.t8 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X364 a_n9707_9395# a_n9329_1995# avss.t304 sky130_fd_pr__res_xhigh_po_1p41 l=35
X365 dvss.t166 sky130_fd_sc_hd__inv_4_0.Y ovout.t9 dvss.t165 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X366 rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.otrip_decoded_avdd[2] avdd.t279 avdd.t278 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X367 comparator_0.vpp comparator_0.vpp avdd.t27 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X368 avdd.t228 comparator_0.vnn comparator_0.vpp avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X369 a_n24817_n11914# a_n24439_n15834# avss.t178 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X370 rstring_mux_0.vtop.t11 rstring_mux_0.ena_b avdd.t406 avdd.t405 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X371 rstring_mux_0.vtrip5.t5 rstring_mux_0.vtrip6.t3 avss.t351 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X372 a_n7751_n3946# a_n8119_n2964# dvss.t305 dvss.t304 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X373 a_9570_n2256# a_9145_n2212# dvss.t73 dvss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X374 a_n20281_n11914# a_n19903_n15834# avss.t243 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X375 dvss.t260 a_10515_n2156# a_10874_n2222# dvss.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X376 avdd.t138 avdd.t136 avdd.t138 avdd.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X377 avdd.t3 a_n3795_n2876# a_n2588_n3212# avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X378 comparator_0.vnn comparator_0.vnn avdd.t227 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X379 schmitt_trigger_0.m.t4 schmitt_trigger_0.in.t5 dvdd.t19 dvdd.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X380 a_7458_n2256# a_7033_n2212# dvss.t245 dvss.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X381 a_n9697_n11914# a_n9319_n15834# avss.t378 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X382 rstring_mux_0.vtrip7.t0 rstring_mux_0.vtrip6.t2 avss.t255 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X383 comparator_0.vn comparator_0.vn avss.t189 avss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X384 dvss.t535 a_n1783_n1230# a_n1683_n1142# dvss.t534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X385 dvss.t293 a_4653_n1142# a_5860_n1478# dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X386 avdd.t306 a_n3102_n3990# a_n3795_n2876# avdd.t305 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X387 comparator_0.vt vbg_1v2.t9 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X388 rstring_mux_0.vtrip15.t4 rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y vin.t91 avdd.t441 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X389 avdd.t374 a_n1683_n1142# a_n990_n2256# avdd.t373 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X390 a_n1683_n2876# a_n1783_n2964# dvss.t397 dvss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X391 ibias_gen_0.ena_b ibias_gen_0.ena avdd.t337 avdd.t336 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X392 a_n3102_n2256# a_n3527_n2212# dvss.t23 dvss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X393 avdd.t135 avdd.t133 avdd.t134 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=8
X394 avss.t118 avss.t117 avss.t118 avss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X395 a_2541_n1142# a_2441_n1230# dvss.t266 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X396 ibias_gen_0.isrc_sel a_10084_n1478# avdd.t355 avdd.t354 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X397 dvss.t439 otrip_decoded[13].t0 a_4553_n1230# dvss.t438 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X398 a_10515_n1026# dcomp avdd.t297 avdd.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X399 avdd.t9 a_n5907_n2876# a_n4700_n3212# avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X400 ibias_gen_0.vn0.t10 vbg_1v2.t10 ibias_gen_0.vstart.t7 avss.t169 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X401 a_9570_n2256# a_9145_n2212# dvss.t71 dvss.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X402 rstring_mux_0.otrip_decoded_avdd[13] a_5860_n1478# dvss.t75 dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X403 dvss.t21 a_n3527_n2212# a_n3102_n2256# dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X404 dvss.t11 a_n1415_n2212# a_n990_n2256# dvss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X405 a_4921_n2212# a_4553_n1230# dvss.t518 dvss.t517 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X406 a_n4405_n11914# a_n4783_n15834# avss.t244 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X407 dvss.t138 a_n3895_n1230# a_n3795_n1142# dvss.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X408 rstring_mux_0.vtop.t0 a_n28219_n15834# avss.t20 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X409 rstring_mux_0.vtop.t10 rstring_mux_0.ena_b avdd.t404 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X410 a_n3795_n2876# a_n3895_n2964# dvss.t233 dvss.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X411 a_n5214_n2256# a_n5639_n2212# dvss.t35 dvss.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X412 rstring_mux_0.otrip_decoded_avdd[12] a_5860_n3212# avdd.t209 avdd.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X413 dvss.t106 otrip_decoded[15].t0 a_6665_n1230# dvss.t105 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X414 comparator_0.vt vbg_1v2.t11 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X415 a_4653_n1142# a_4553_n1230# dvss.t516 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X416 a_n990_n2256# a_n1415_n2212# dvss.t9 dvss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X417 a_n1415_n2212# a_n1783_n1230# dvdd.t143 dvdd.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X418 dvss.t512 a_n6007_n2964# a_n5907_n2876# dvss.t511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X419 dvss.t409 a_4553_n2964# a_4653_n2876# dvss.t408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X420 avdd.t315 a_n8019_n2876# a_n6812_n3212# avdd.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X421 ibias_gen_0.vp1.t3 ibias_gen_0.isrc_sel ibias_gen_0.vp.t3 avss.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X422 a_n23305_n11914# a_n22927_n15834# avss.t338 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X423 ibias_gen_0.vstart.t6 vbg_1v2.t12 ibias_gen_0.vn0.t11 avss.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X424 ovout.t8 sky130_fd_sc_hd__inv_4_0.Y dvss.t164 dvss.t163 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X425 dvss.t89 a_6665_n1230# a_6765_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X426 rstring_mux_0.otrip_decoded_avdd[15] a_7972_n1478# dvss.t458 dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X427 dvss.t33 a_n5639_n2212# a_n5214_n2256# dvss.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X428 rstring_mux_0.vtop.t9 rstring_mux_0.ena_b avdd.t402 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X429 a_n23305_n11914# a_n23683_n15834# avss.t54 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X430 a_n5907_n2876# a_n6007_n2964# dvss.t510 dvss.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X431 dvdd.t93 otrip_decoded[10].t1 a_2441_n2964# dvdd.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X432 ibias_gen_0.isrc_sel_b avdd.t131 ibias_gen_0.ena_b avdd.t132 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X433 dvdd.t3 isrc_sel.t1 a_8777_n1230# dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X434 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t9 dvss.t347 dvss.t346 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X435 a_n7326_n2256# a_n7751_n2212# dvss.t61 dvss.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X436 a_n8185_n11914# a_n7807_n15834# avss.t328 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X437 vin.t57 rstring_mux_0.otrip_decoded_b_avdd[8] rstring_mux_0.vtrip8.t5 avdd.t349 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X438 avdd.t194 a_429_n2876# a_1636_n3212# avdd.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X439 comparator_0.vt avss.t388 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X440 a_n23050_n2937# a_n22672_n10337# avss.t199 sky130_fd_pr__res_xhigh_po_1p41 l=35
X441 a_6765_n1142# a_6665_n1230# dvss.t88 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X442 a_n3527_n2212# a_n3895_n1230# dvdd.t27 dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X443 comparator_0.ena_b ibias_gen_0.ena avss.t322 avss.t321 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X444 dvss.t303 a_n8119_n2964# a_n8019_n2876# dvss.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X445 a_n11209_n11914# a_n11587_n15834# avss.t311 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X446 dvss.t425 a_6665_n2964# a_6765_n2876# dvss.t424 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X447 a_n13487_9395# a_n13865_1995# avss.t281 sky130_fd_pr__res_xhigh_po_1p41 l=35
X448 comparator_0.vnn avss.t389 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X449 a_1122_n2256# a_697_n2212# dvss.t279 dvss.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X450 a_n22294_n2937# a_n21916_n10337# avss.t204 sky130_fd_pr__res_xhigh_po_1p41 l=35
X451 dvss.t80 a_8777_n1230# a_8877_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X452 dvss.t59 a_n7751_n2212# a_n7326_n2256# dvss.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X453 rstring_mux_0.vtrip4.t5 rstring_mux_0.otrip_decoded_b_avdd[4] vin.t90 avdd.t440 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X454 dvss.t292 a_697_n3946# a_1122_n3990# dvss.t291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X455 vin.t15 rstring_mux_0.otrip_decoded_b_avdd[12] rstring_mux_0.vtrip12.t1 avdd.t212 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X456 a_8877_n2876# a_8777_n2964# dvss.t331 dvss.t330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X457 avdd.t245 comparator_0.n0 comparator_0.n1 avdd.t244 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X458 avdd.t359 a_8877_n1142# a_9570_n2256# avdd.t358 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X459 vin.t35 avss.t115 vin.t35 avss.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X460 avdd.t184 a_1122_n3990# a_429_n2876# avdd.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X461 avdd.t26 comparator_0.vpp comparator_0.vpp avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X462 schmitt_trigger_0.out.t2 schmitt_trigger_0.m.t16 dvdd.t107 dvdd.t106 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X463 a_429_n2876# a_329_n2964# dvss.t192 dvss.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X464 a_8877_n1142# a_8777_n1230# dvss.t79 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X465 a_n5639_n2212# a_n6007_n1230# dvdd.t135 dvdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X466 dvss.t329 a_8777_n2964# a_8877_n2876# dvss.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X467 dvdd.t43 sky130_fd_sc_hd__inv_4_0.Y ovout.t23 dvdd.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X468 a_n27085_n11914# a_n26707_n15834# avss.t205 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X469 rstring_mux_0.vtop.t8 rstring_mux_0.ena_b avdd.t400 avdd.t399 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X470 a_3234_n2256# a_2809_n2212# dvss.t373 dvss.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X471 rstring_mux_0.otrip_decoded_b_avdd[9] rstring_mux_0.otrip_decoded_avdd[9] avdd.t265 avdd.t264 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X472 a_n11219_9395# a_n10841_1995# avss.t332 sky130_fd_pr__res_xhigh_po_1p41 l=35
X473 dvss.t190 a_329_n2964# a_429_n2876# dvss.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X474 comparator_0.vnn vbg_1v2.t13 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X475 avdd.t398 rstring_mux_0.ena_b rstring_mux_0.vtop.t7 avdd.t397 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X476 a_8877_n2876# a_8777_n2964# dvss.t327 dvss.t326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X477 avdd.t130 avdd.t128 avdd.t129 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=8
X478 ibias_gen_0.vp0.t9 ibias_gen_0.ena avdd.t335 avdd.t334 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X479 vin.t78 avdd.t126 vin.t78 avdd.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X480 rstring_mux_0.otrip_decoded_b_avdd[9] rstring_mux_0.otrip_decoded_avdd[9] avss.t223 avss.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X481 rstring_mux_0.otrip_decoded_b_avdd[13] rstring_mux_0.otrip_decoded_avdd[13] avdd.t430 avdd.t429 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X482 avdd.t371 a_3234_n3990# a_2541_n2876# avdd.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X483 avdd.t250 a_6765_n2876# a_7972_n3212# avdd.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X484 rstring_mux_0.otrip_decoded_avdd[8] a_1636_n3212# avdd.t210 avdd.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X485 a_5346_n3990# a_4921_n3946# dvss.t221 dvss.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X486 ibias_gen_0.vn0.t0 ibias_gen_0.ena_b avss.t3 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X487 dvss.t455 a_6765_n1142# a_7972_n1478# dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X488 dvdd.t95 otrip_decoded[8].t1 a_329_n2964# dvdd.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X489 a_10515_n2156# a_10515_n1026# avdd.t298 avdd.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X490 rstring_mux_0.vtop.t6 rstring_mux_0.ena_b avdd.t396 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X491 comparator_0.vt vin.t101 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X492 vin.t88 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.vtrip1.t4 avss.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X493 comparator_0.vpp comparator_0.vnn avdd.t226 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X494 avdd.t25 comparator_0.vpp comparator_0.vnn avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X495 a_n9707_9395# a_n10085_1995# avss.t330 sky130_fd_pr__res_xhigh_po_1p41 l=35
X496 avdd.t326 a_n5907_n1142# a_n5214_n2256# avdd.t325 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X497 dvss.t533 a_n1783_n1230# a_n1683_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X498 avdd.t225 comparator_0.vnn comparator_0.vm avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X499 avss.t114 avss.t113 ibias_gen_0.ve.t3 avss sky130_fd_pr__pnp_05v5_W0p68L0p68
**devattr s=18496,544 d=4547244,10712
X500 dvdd.t124 otrip_decoded[13].t1 a_4553_n1230# dvdd.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X501 rstring_mux_0.otrip_decoded_avdd[10] a_3748_n3212# avdd.t281 avdd.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X502 schmitt_trigger_0.in.t6 dvss.t115 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X503 a_7458_n3990# a_7033_n3946# dvss.t130 dvss.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X504 avdd.t293 a_5346_n3990# a_4653_n2876# avdd.t292 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X505 a_7691_n11914# a_7313_n15834# avss.t242 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X506 vin.t77 avdd.t124 vin.t77 avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X507 rstring_mux_0.otrip_decoded_b_avdd[3] rstring_mux_0.otrip_decoded_avdd[3] avss.t9 avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X508 avss.t249 comparator_0.vm comparator_0.n0 avss.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X509 avss.t112 avss.t110 avss.t111 avss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X510 a_n1683_n1142# a_n1783_n1230# dvss.t532 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X511 vin.t34 avss.t108 vin.t34 avss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X512 comparator_0.vnn vbg_1v2.t14 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X513 a_4921_n2212# a_4553_n1230# dvdd.t141 dvdd.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X514 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t10 dvss.t349 dvss.t348 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X515 a_9570_n2256# a_9145_n2212# dvss.t69 dvss.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X516 comparator_0.vnn avss.t390 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X517 dvss.t265 a_2441_n1230# a_2541_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X518 dvss.t7 a_n1415_n2212# a_n990_n2256# dvss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X519 schmitt_trigger_0.in.t7 dvss.t116 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X520 ibias_gen_0.vn1.t2 avss.t106 ibias_gen_0.vp1.t1 avss.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X521 avdd.t382 a_n8019_n1142# a_n7326_n2256# avdd.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X522 dvss.t136 a_n3895_n1230# a_n3795_n1142# dvss.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X523 a_2541_n2876# a_2441_n2964# dvss.t341 dvss.t340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X524 vin.t25 rstring_mux_0.otrip_decoded_avdd[14] rstring_mux_0.vtrip14.t3 avss.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X525 a_n990_n3990# a_n1415_n3946# dvss.t361 dvss.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X526 ibias_gen_0.vn0.t12 vbg_1v2.t15 ibias_gen_0.vstart.t5 avss.t171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X527 dvdd.t99 otrip_decoded[15].t1 a_6665_n1230# dvdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X528 a_n3795_n2876# a_n3895_n2964# dvss.t231 dvss.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X529 dvss.t387 a_n5907_n1142# a_n4700_n1478# dvss.t386 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X530 a_n5214_n2256# a_n5639_n2212# dvss.t31 dvss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X531 avdd.t308 a_7458_n3990# a_6765_n2876# avdd.t307 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X532 a_n7751_n3946# a_n8119_n2964# dvdd.t85 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X533 dvss.t162 sky130_fd_sc_hd__inv_4_0.Y ovout.t7 dvss.t161 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X534 a_n3102_n2256# a_n3527_n2212# dvss.t19 dvss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X535 a_n990_n2256# a_n1415_n2212# dvss.t5 dvss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X536 dvss.t476 a_10874_n2222# vl.t1 dvss.t475 sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X537 comparator_0.vpp comparator_0.vnn avdd.t224 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X538 vin.t61 rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.vtrip2.t2 avdd.t375 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X539 rstring_mux_0.otrip_decoded_avdd[9] a_1636_n1478# dvss.t431 dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X540 dvss.t339 a_2441_n2964# a_2541_n2876# dvss.t338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X541 rstring_mux_0.vtrip8.t4 rstring_mux_0.otrip_decoded_b_avdd[8] vin.t58 avdd.t348 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X542 rstring_mux_0.vtrip0.t1 rstring_mux_0.otrip_decoded_b_avdd[0] vin.t20 avdd.t263 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X543 dvss.t488 a_n6007_n1230# a_n5907_n1142# dvss.t487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X544 rstring_mux_0.vtrip15.t1 rstring_mux_0.otrip_decoded_avdd[15] vin.t11 avss.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X545 comparator_0.n0 comparator_0.ena_b avss.t182 avss.t181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X546 a_n5907_n2876# a_n6007_n2964# dvss.t508 dvss.t507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X547 a_n5907_n2876# a_n6007_n2964# dvss.t506 dvss.t505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X548 a_4653_n2876# a_4553_n2964# dvss.t407 dvss.t406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X549 avss.t343 rstring_mux_0.ena_b rstring_mux_0.vtop.t17 avss.t342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X550 avdd.t289 a_2541_n2876# a_3748_n3212# avdd.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X551 avss.t33 comparator_0.n1 dcomp avss.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X552 avss.t292 ibias_gen_0.vn1.t15 ibias_gen_0.vp1.t9 avss.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X553 a_n7326_n2256# a_n7751_n2212# dvss.t57 dvss.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X554 vin.t0 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.vtrip3.t0 avss.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X555 rstring_mux_0.vtrip12.t0 rstring_mux_0.otrip_decoded_b_avdd[12] vin.t14 avdd.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X556 avdd.t256 a_9570_n3990# a_8877_n2876# avdd.t255 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X557 a_n8019_n1142# a_n8119_n1230# dvss.t94 dvss.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X558 a_n1415_n3946# a_n1783_n2964# dvss.t395 dvss.t394 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X559 ibias_gen_0.vstart.t4 vbg_1v2.t16 ibias_gen_0.vn0.t13 avss.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X560 dvss.t301 a_n8119_n2964# a_n8019_n2876# dvss.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X561 a_n8185_n11914# a_n8563_n15834# avss.t312 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X562 vin.t33 avss.t104 vin.t33 avss.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X563 vin.t16 rstring_mux_0.otrip_decoded_avdd[6] rstring_mux_0.vtrip6.t1 avss.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X564 a_1122_n2256# a_697_n2212# dvss.t277 dvss.t276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X565 comparator_0.vt avss.t391 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X566 avss.t103 avss.t101 avss.t102 avss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X567 dvdd.t41 sky130_fd_sc_hd__inv_4_0.Y ovout.t22 dvdd.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X568 a_10874_n1026# a_10515_n1026# dvss.t315 dvss.t312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X569 a_n8019_n2876# a_n8119_n2964# dvss.t299 dvss.t298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X570 dvss.t474 ena.t0 a_8777_n2964# dvss.t473 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X571 a_6765_n2876# a_6665_n2964# dvss.t423 dvss.t422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X572 avdd.t123 avdd.t121 avdd.t123 avdd.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X573 dvss.t371 a_2809_n2212# a_3234_n2256# dvss.t370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X574 a_n8019_n2876# a_n8119_n2964# dvss.t297 dvss.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X575 rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.otrip_decoded_avdd[0] avdd.t420 avdd.t419 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X576 avdd.t257 a_4653_n2876# a_5860_n3212# avdd.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X577 dvss.t309 dcomp a_10515_n1026# dvss.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X578 dvss.t275 a_697_n2212# a_1122_n2256# dvss.t274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X579 rstring_mux_0.vtrip1.t2 rstring_mux_0.vtrip0.t3 avss.t313 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X580 a_n3527_n3946# a_n3895_n2964# dvss.t229 dvss.t228 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X581 a_429_n2876# a_329_n2964# dvss.t188 dvss.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X582 vin.t38 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.vtrip7.t1 avss.t266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X583 avdd.t120 avdd.t118 avdd.t119 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=8
X584 avdd.t117 avdd.t116 avdd.t117 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=8
X585 a_n3649_n11914# rstring_mux_0.vtrip0.t2 avss.t302 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X586 avdd.t223 comparator_0.vnn comparator_0.vnn avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X587 a_n14243_9395# a_n13865_1995# avss.t272 sky130_fd_pr__res_xhigh_po_1p41 l=35
X588 vin.t26 rstring_mux_0.otrip_decoded_avdd[12] rstring_mux_0.vtrip12.t3 avss.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X589 dvss.t351 schmitt_trigger_0.out.t11 sky130_fd_sc_hd__inv_4_0.Y dvss.t350 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X590 a_3234_n2256# a_2809_n2212# dvss.t369 dvss.t368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X591 a_n27085_n11914# a_n27463_n15834# avss.t273 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X592 avdd.t352 a_n3795_n1142# a_n3102_n2256# avdd.t351 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X593 dvss.t204 a_2809_n3946# a_3234_n3990# dvss.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X594 dvdd.t39 sky130_fd_sc_hd__inv_4_0.Y ovout.t21 dvdd.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X595 ovout.t6 sky130_fd_sc_hd__inv_4_0.Y dvss.t160 dvss.t159 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X596 dvss.t186 a_329_n2964# a_429_n2876# dvss.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X597 rstring_mux_0.otrip_decoded_avdd[7] a_n476_n1478# dvss.t282 dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X598 avss.t100 avss.t99 avss.t100 avss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X599 dvss.t468 a_4921_n2212# a_5346_n2256# dvss.t467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X600 vin.t10 rstring_mux_0.otrip_decoded_avdd[15] rstring_mux_0.vtrip15.t0 avss.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X601 comparator_0.vt avss.t392 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X602 avss.t356 a_n27208_n10337# avss.t355 sky130_fd_pr__res_xhigh_po_1p41 l=35
X603 a_n5639_n3946# a_n6007_n2964# dvss.t504 dvss.t503 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X604 a_n21793_n11914# a_n22171_n15834# avss.t377 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X605 rstring_mux_0.vtrip13.t4 rstring_mux_0.otrip_decoded_avdd[13] vin.t79 avss.t364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X606 comparator_0.vnn avss.t393 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X607 ibias_gen_0.ibias ibias_gen_0.vp.t10 avdd.t51 avdd.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X608 rstring_mux_0.vtrip5.t3 rstring_mux_0.otrip_decoded_b_avdd[5] vin.t54 avdd.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X609 a_5346_n2256# a_4921_n2212# dvss.t466 dvss.t465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X610 a_n22549_n11914# a_n22171_n15834# avss.t24 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X611 rstring_mux_0.otrip_decoded_b_avdd[11] rstring_mux_0.otrip_decoded_avdd[11] avdd.t432 avdd.t431 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X612 vin.t18 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.vtrip5.t0 avss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X613 comparator_0.vt vin.t102 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X614 rstring_mux_0.vtrip15.t2 rstring_mux_0.vtrip14.t1 avss.t165 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X615 a_9570_n3990# a_9145_n3946# dvss.t43 dvss.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X616 avdd.t273 a_429_n1142# a_1122_n2256# avdd.t272 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X617 a_n6673_n11914# a_n7051_n15834# avss.t55 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X618 avdd.t115 avdd.t113 avdd.t114 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=8
X619 dvss.t243 a_7033_n2212# a_7458_n2256# dvss.t242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X620 a_n15479_n3901# ibias_gen_0.isrc_sel ibias_gen_0.vn1.t3 avss.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X621 dvss.t384 a_2541_n1142# a_3748_n1478# dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X622 rstring_mux_0.otrip_decoded_avdd[2] a_n4700_n3212# dvss.t472 dvss.t471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X623 a_n10453_n11914# a_n10075_n15834# avss.t58 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X624 a_n7429_n11914# a_n7051_n15834# avss.t152 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X625 rstring_mux_0.otrip_decoded_b_avdd[11] rstring_mux_0.otrip_decoded_avdd[11] avss.t368 avss.t367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X626 a_7458_n3990# a_7033_n3946# dvss.t128 dvss.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X627 ovout.t5 sky130_fd_sc_hd__inv_4_0.Y dvss.t158 dvss.t157 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X628 dvss.t393 a_n1783_n2964# a_n1683_n2876# dvss.t392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X629 ibias_gen_0.vp0.t0 ibias_gen_0.vn0.t20 ibias_gen_0.vr.t0 avss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X630 comparator_0.vpp comparator_0.vpp avdd.t24 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X631 comparator_0.vnn comparator_0.vpp avdd.t23 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X632 a_2809_n2212# a_2441_n1230# dvss.t264 dvss.t263 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X633 dvss.t17 a_n3527_n2212# a_n3102_n2256# dvss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X634 avdd.t192 a_n5214_n3990# a_n5907_n2876# avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X635 avdd.t22 comparator_0.vpp comparator_0.vpp avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X636 comparator_0.vnn vbg_1v2.t17 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X637 a_n3102_n3990# a_n3527_n3946# dvss.t449 dvss.t448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X638 dvdd.t21 schmitt_trigger_0.in.t8 schmitt_trigger_0.m.t5 dvdd.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X639 a_2541_n2876# a_2441_n2964# dvss.t337 dvss.t336 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X640 rstring_mux_0.otrip_decoded_b_avdd[5] rstring_mux_0.otrip_decoded_avdd[5] avdd.t239 avdd.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X641 dvss.t415 otrip_decoded[12].t0 a_4553_n2964# dvss.t414 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X642 avss.t98 avss.t95 avss.t97 avss.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X643 comparator_0.vnn avss.t394 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X644 avdd.t317 a_2541_n1142# a_3234_n2256# avdd.t316 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X645 dvss.t67 a_9145_n2212# a_9570_n2256# dvss.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X646 rstring_mux_0.vtrip7.t5 rstring_mux_0.otrip_decoded_b_avdd[7] vin.t60 avdd.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X647 dvdd.t37 sky130_fd_sc_hd__inv_4_0.Y ovout.t20 dvdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X648 a_n25573_n11914# a_n25951_n15834# avss.t370 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X649 vin.t2 rstring_mux_0.otrip_decoded_avdd[10] rstring_mux_0.vtrip10.t0 avss.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X650 comparator_0.n0 comparator_0.vm avss.t248 avss.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X651 a_n3102_n2256# a_n3527_n2212# dvss.t15 dvss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X652 rstring_mux_0.otrip_decoded_avdd[0] a_n6812_n3212# dvss.t253 dvss.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X653 a_9570_n3990# a_9145_n3946# dvss.t41 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X654 a_4921_n3946# a_4553_n2964# dvss.t405 dvss.t404 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X655 dvss.t359 a_n1415_n3946# a_n990_n3990# dvss.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X656 dvss.t447 a_n3527_n3946# a_n3102_n3990# dvss.t446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X657 comparator_0.vt vin.t103 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X658 dvss.t227 a_n3895_n2964# a_n3795_n2876# dvss.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X659 vin.t76 avdd.t111 vin.t76 avdd.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X660 rstring_mux_0.otrip_decoded_b_avdd[10] rstring_mux_0.otrip_decoded_avdd[10] avdd.t39 avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X661 a_7033_n2212# a_6665_n1230# dvss.t87 dvss.t86 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X662 avss.t210 comparator_0.n0 comparator_0.n1 avss.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X663 dvss.t29 a_n5639_n2212# a_n5214_n2256# dvss.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X664 a_6179_n11914# a_5801_n15834# avss.t216 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X665 avdd.t277 a_n7326_n3990# a_n8019_n2876# avdd.t276 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X666 dvss.t515 a_4553_n1230# a_4653_n1142# dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X667 a_n13477_n11914# a_n13855_n15834# avss.t310 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X668 a_n5214_n3990# a_n5639_n3946# dvss.t531 dvss.t530 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X669 dvss.t413 otrip_decoded[7].t0 a_n1783_n1230# dvss.t412 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X670 dvss.t251 otrip_decoded[14].t0 a_6665_n2964# dvss.t250 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X671 avdd.t287 a_4653_n1142# a_5346_n2256# avdd.t286 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X672 vin.t89 rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.vtrip4.t4 avdd.t439 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X673 a_n990_n3990# a_n1415_n3946# dvss.t357 dvss.t356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X674 a_4653_n2876# a_4553_n2964# dvss.t403 dvss.t402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X675 avdd.t110 avdd.t109 avdd.t110 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=8
X676 dvdd.t35 sky130_fd_sc_hd__inv_4_0.Y ovout.t19 dvdd.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X677 vin.t84 rstring_mux_0.otrip_decoded_b_avdd[14] rstring_mux_0.vtrip14.t5 avdd.t434 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X678 avdd.t20 comparator_0.vpp comparator_0.vnn avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X679 avdd.t59 comparator_0.n1 dcomp avdd.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X680 a_n5214_n2256# a_n5639_n2212# dvss.t27 dvss.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X681 dcomp comparator_0.n1 avdd.t57 avdd.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X682 comparator_0.vm comparator_0.vnn avdd.t222 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X683 dvss.t529 a_n5639_n3946# a_n5214_n3990# dvss.t528 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X684 dvss.t421 a_6665_n2964# a_6765_n2876# dvss.t420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X685 rstring_mux_0.otrip_decoded_b_avdd[7] rstring_mux_0.otrip_decoded_avdd[7] avdd.t300 avdd.t299 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X686 comparator_0.vnn avss.t395 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X687 avss.t31 comparator_0.n1 dcomp avss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X688 a_1122_n2256# a_697_n2212# dvss.t273 dvss.t272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X689 a_9145_n2212# a_8777_n1230# dvss.t77 dvss.t76 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X690 dvss.t55 a_n7751_n2212# a_n7326_n2256# dvss.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X691 rstring_mux_0.vtrip11.t1 rstring_mux_0.vtrip12.t2 avss.t217 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X692 a_n7326_n3990# a_n7751_n3946# dvss.t484 dvss.t483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X693 dvss.t454 otrip_decoded[5].t0 a_n3895_n1230# dvss.t453 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X694 avdd.t378 a_6765_n1142# a_7458_n2256# avdd.t377 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X695 a_6765_n2876# a_6665_n2964# dvss.t419 dvss.t418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X696 dvdd.t122 dvdd.t120 schmitt_trigger_0.m.t13 dvdd.t121 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X697 a_697_n2212# a_329_n1230# dvss.t209 dvss.t208 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X698 ovout.t4 sky130_fd_sc_hd__inv_4_0.Y dvss.t156 dvss.t155 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X699 a_n17257_n11914# a_n16879_n15834# avss.t18 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X700 a_1122_n3990# a_697_n3946# dvss.t290 dvss.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X701 a_n26074_n2937# a_n25696_n10337# avss.t319 sky130_fd_pr__res_xhigh_po_1p41 l=35
X702 dvss.t482 a_n7751_n3946# a_n7326_n3990# dvss.t481 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X703 dvss.t325 a_8777_n2964# a_8877_n2876# dvss.t324 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X704 a_n11219_9395# a_n11597_1995# avss.t214 sky130_fd_pr__res_xhigh_po_1p41 l=35
X705 a_n17257_n11914# a_n17635_n15834# avss.t215 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X706 rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y rstring_mux_0.otrip_decoded_avdd[15] avdd.t186 avdd.t185 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X707 a_n12731_9395# a_n12353_1995# avss.t254 sky130_fd_pr__res_xhigh_po_1p41 l=35
X708 a_429_n1142# a_329_n1230# dvss.t207 dvss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X709 a_3234_n2256# a_2809_n2212# dvss.t367 dvss.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X710 a_n25318_n2937# a_n24940_n10337# avss.t352 sky130_fd_pr__res_xhigh_po_1p41 l=35
X711 avdd.t243 a_8877_n2876# a_10084_n3212# avdd.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X712 vin.t53 rstring_mux_0.otrip_decoded_b_avdd[5] rstring_mux_0.vtrip5.t2 avdd.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X713 rstring_mux_0.otrip_decoded_avdd[14] a_7972_n3212# dvss.t49 dvss.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X714 comparator_0.vnn vbg_1v2.t18 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X715 dvss.t452 otrip_decoded[3].t0 a_n6007_n1230# dvss.t451 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X716 a_8877_n2876# a_8777_n2964# dvss.t323 dvss.t322 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X717 avss.t162 ibias_gen_0.isrc_sel ibias_gen_0.vn0.t6 avss.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X718 dvss.t464 a_4921_n2212# a_5346_n2256# dvss.t463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X719 avss.t160 ibias_gen_0.isrc_sel ibias_gen_0.isrc_sel_b avss.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X720 ovout.t3 sky130_fd_sc_hd__inv_4_0.Y dvss.t154 dvss.t153 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X721 a_10715_n11914# a_10337_n15834# avss.t300 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X722 a_n1415_n3946# a_n1783_n2964# dvdd.t109 dvdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X723 a_n11965_n11914# a_n12343_n15834# avss.t316 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X724 a_n8941_n11914# a_n9319_n15834# avss.t317 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X725 a_4667_n11914# a_4289_n15834# avss.t318 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X726 a_3234_n3990# a_2809_n3946# dvss.t202 dvss.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X727 comparator_0.vnn comparator_0.vnn avdd.t221 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X728 comparator_0.vt avss.t396 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X729 a_n12721_n11914# a_n12343_n15834# avss.t353 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X730 a_4667_n11914# a_5045_n15834# avss.t354 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X731 a_n22294_n2937# a_n22672_n10337# avss.t315 sky130_fd_pr__res_xhigh_po_1p41 l=35
X732 dvdd.t65 schmitt_trigger_0.out.t12 schmitt_trigger_0.m.t10 dvdd.t64 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X733 a_5346_n2256# a_4921_n2212# dvss.t462 dvss.t461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X734 ibias_gen_0.vp1.t17 ibias_gen_0.isrc_sel_b ibias_gen_0.vp.t6 avdd.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X735 avdd.t394 rstring_mux_0.ena_b rstring_mux_0.vtop.t5 avdd.t393 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X736 dvss.t108 otrip_decoded[1].t0 a_n8119_n1230# dvss.t107 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X737 dvdd.t97 ena.t1 a_8777_n2964# dvdd.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X738 a_n24562_n2937# a_n24940_n10337# avss.t252 sky130_fd_pr__res_xhigh_po_1p41 l=35
X739 a_n21538_n2937# a_n21916_n10337# avss.t253 sky130_fd_pr__res_xhigh_po_1p41 l=35
X740 dvss.t241 a_7033_n2212# a_7458_n2256# dvss.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X741 a_n3527_n3946# a_n3895_n2964# dvdd.t79 dvdd.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X742 ibias_gen_0.vstart.t3 vbg_1v2.t19 ibias_gen_0.vn0.t14 avss.t173 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X743 avss.t284 ibias_gen_0.vn1.t4 ibias_gen_0.vn1.t5 avss.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X744 rstring_mux_0.otrip_decoded_avdd[6] a_n476_n3212# dvss.t47 dvss.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X745 avdd.t75 a_n1683_n2876# a_n990_n3990# avdd.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X746 vin.t59 rstring_mux_0.otrip_decoded_b_avdd[7] rstring_mux_0.vtrip7.t4 avdd.t356 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X747 a_n23806_n2937# a_n24184_n10337# avss.t381 sky130_fd_pr__res_xhigh_po_1p41 l=35
X748 avss.t1 ibias_gen_0.ena_b ibias_gen_0.vn1.t0 avss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X749 a_2809_n2212# a_2441_n1230# dvdd.t83 dvdd.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X750 dvss.t391 a_n1783_n2964# a_n1683_n2876# dvss.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X751 a_n27841_n11914# a_n28219_n15834# avss.t230 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X752 a_7458_n2256# a_7033_n2212# dvss.t239 dvss.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X753 avdd.t392 rstring_mux_0.ena_b rstring_mux_0.vtop.t4 avdd.t391 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X754 ibias_gen_0.ena a_10084_n3212# avdd.t417 avdd.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X755 rstring_mux_0.otrip_decoded_b_avdd[13] rstring_mux_0.otrip_decoded_avdd[13] avss.t363 avss.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X756 comparator_0.vpp vin.t104 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X757 avdd.t108 avdd.t106 avdd.t107 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=8
X758 avdd.t105 avdd.t104 avdd.t105 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=8
X759 vin.t21 rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.vtrip0.t0 avdd.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X760 ibias_gen_0.isrc_sel a_10084_n1478# dvss.t434 dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X761 avss.t94 avss.t93 avss.t94 avss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X762 dvss.t65 a_9145_n2212# a_9570_n2256# dvss.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X763 a_n1683_n2876# a_n1783_n2964# dvss.t389 dvss.t388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X764 a_n15745_n11914# a_n16123_n15834# avss.t295 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X765 a_8447_n11914# a_8069_n15834# avss.t296 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X766 ibias_gen_0.ve.t2 avss.t90 avss.t92 avss.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X767 rstring_mux_0.otrip_decoded_avdd[3] a_n4700_n1478# avdd.t182 avdd.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X768 a_n5639_n3946# a_n6007_n2964# dvdd.t137 dvdd.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X769 a_9570_n3990# a_9145_n3946# dvss.t39 dvss.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X770 a_n16501_n11914# a_n16123_n15834# avss.t299 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X771 a_7033_n2212# a_6665_n1230# dvdd.t9 dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X772 dvss.t335 a_2441_n2964# a_2541_n2876# dvss.t334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X773 dvss.t355 a_n1415_n3946# a_n990_n3990# dvss.t354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X774 avdd.t19 comparator_0.vpp comparator_0.vnn avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X775 dvdd.t33 sky130_fd_sc_hd__inv_4_0.Y ovout.t18 dvdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X776 ovout.t2 sky130_fd_sc_hd__inv_4_0.Y dvss.t152 dvss.t151 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X777 dvss.t225 a_n3895_n2964# a_n3795_n2876# dvss.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X778 rstring_mux_0.vtrip14.t4 rstring_mux_0.otrip_decoded_b_avdd[14] vin.t83 avdd.t433 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X779 ibias_gen_0.vp1.t10 ibias_gen_0.vn1.t16 avss.t293 avss.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X780 dvss.t433 a_n3795_n1142# a_n2588_n1478# dvss.t432 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X781 avss.t294 ibias_gen_0.vn1.t17 ibias_gen_0.vp1.t11 avss.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X782 dvdd.t115 otrip_decoded[7].t1 a_n1783_n1230# dvdd.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X783 comparator_0.vt vin.t105 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X784 a_n20782_n2937# a_n20404_n10337# avss.t17 sky130_fd_pr__res_xhigh_po_1p41 l=35
X785 dvss.t258 a_10515_n2156# a_10874_n2222# dvss.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X786 a_n5214_n3990# a_n5639_n3946# dvss.t527 dvss.t526 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X787 dcomp comparator_0.n1 avdd.t55 avdd.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X788 vin.t32 avdd.t102 vin.t32 avdd.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X789 a_n990_n3990# a_n1415_n3946# dvss.t353 dvss.t352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X790 a_n3102_n3990# a_n3527_n3946# dvss.t445 dvss.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X791 a_3155_n11914# a_3533_n15834# avss.t265 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X792 rstring_mux_0.vtrip1.t3 rstring_mux_0.otrip_decoded_avdd[1] vin.t87 avss.t371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X793 rstring_mux_0.otrip_decoded_avdd[1] a_n6812_n1478# avdd.t207 avdd.t206 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X794 a_n11209_n11914# a_n10831_n15834# avss.t336 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X795 dvss.t314 a_10515_n1026# a_10874_n1026# dvss.t312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X796 a_n7326_n2256# a_n7751_n2212# dvss.t53 dvss.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X797 dvss.t51 a_n1683_n2876# a_n476_n3212# dvss.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X798 a_10874_n2222# a_10515_n2156# dvss.t256 dvss.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X799 avdd.t101 avdd.t98 avdd.t100 avdd.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=4
X800 a_9145_n2212# a_8777_n1230# dvdd.t7 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X801 dvss.t502 a_n6007_n2964# a_n5907_n2876# dvss.t501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X802 avdd.t390 rstring_mux_0.ena_b rstring_mux_0.vtop.t3 avdd.t389 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X803 ovout.t1 sky130_fd_sc_hd__inv_4_0.Y dvss.t150 dvss.t149 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X804 avdd.t97 avdd.t95 avdd.t96 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=8
X805 comparator_0.vt avss.t397 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X806 comparator_0.vnn vbg_1v2.t20 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X807 dvdd.t130 otrip_decoded[5].t1 a_n3895_n1230# dvdd.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X808 a_10874_n1026# a_10515_n1026# dvss.t313 dvss.t312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X809 a_n7326_n3990# a_n7751_n3946# dvss.t480 dvss.t479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X810 a_697_n2212# a_329_n1230# dvdd.t77 dvdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X811 a_n8019_n2876# a_n8119_n2964# dvss.t295 dvss.t294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X812 a_n19525_n11914# a_n19903_n15834# avss.t282 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X813 dvdd.t117 otrip_decoded[12].t1 a_4553_n2964# dvdd.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X814 comparator_0.vpp comparator_0.vpp avdd.t18 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X815 comparator_0.vnn comparator_0.vpp avdd.t16 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X816 rstring_mux_0.vtrip7.t3 rstring_mux_0.vtrip8.t3 avss.t279 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X817 vin.t22 rstring_mux_0.otrip_decoded_avdd[9] rstring_mux_0.vtrip9.t0 avss.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X818 a_1122_n3990# a_697_n3946# dvss.t288 dvss.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X819 avdd.t220 comparator_0.vnn comparator_0.vnn avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X820 ibg_200n ibias_gen_0.ena a_n15479_n3901# avss.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X821 avdd.t388 rstring_mux_0.ena_b rstring_mux_0.vtop.t2 avdd.t387 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X822 a_4921_n3946# a_4553_n2964# dvdd.t111 dvdd.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X823 avdd.t241 a_8877_n2876# a_9570_n3990# avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X824 a_n16775_n2223# ibias_gen_0.ena_b ibias_gen_0.vstart.t0 avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X825 vin.t50 rstring_mux_0.otrip_decoded_b_avdd[9] rstring_mux_0.vtrip9.t4 avdd.t310 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X826 avdd.t367 ibias_gen_0.vp0.t12 ibias_gen_0.vn0.t17 avdd.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X827 a_6935_n11914# a_6557_n15834# avss.t261 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X828 dvss.t200 a_2809_n3946# a_3234_n3990# dvss.t199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X829 dvdd.t128 otrip_decoded[3].t1 a_n6007_n1230# dvdd.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X830 a_6935_n11914# a_7313_n15834# avss.t262 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X831 dvss.t286 a_697_n3946# a_1122_n3990# dvss.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X832 ibias_gen_0.ve.t0 ibias_gen_0.vn0.t1 ibias_gen_0.vn0.t2 avss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X833 a_n14989_n11914# a_n14611_n15834# avss.t259 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X834 a_n3649_n11914# a_n4027_n15834# avss.t260 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X835 rstring_mux_0.vtrip3.t4 rstring_mux_0.otrip_decoded_b_avdd[3] vin.t5 avdd.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X836 dvdd.t81 otrip_decoded[14].t1 a_6665_n2964# dvdd.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X837 vin.t13 rstring_mux_0.otrip_decoded_avdd[8] rstring_mux_0.vtrip8.t0 avss.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X838 a_n4405_n11914# a_n4027_n15834# avss.t276 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X839 avss.t187 comparator_0.vn comparator_0.vt avss.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X840 comparator_0.vnn vbg_1v2.t21 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X841 a_3234_n3990# a_2809_n3946# dvss.t198 dvss.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X842 dvdd.t31 sky130_fd_sc_hd__inv_4_0.Y ovout.t17 dvdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X843 a_10715_n11914# avss.t278 avss.t277 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X844 ibias_gen_0.vn0.t15 vbg_1v2.t22 ibias_gen_0.vstart.t2 avss.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X845 rstring_mux_0.otrip_decoded_avdd[15] a_7972_n1478# avdd.t384 avdd.t379 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X846 dvdd.t13 otrip_decoded[1].t1 a_n8119_n1230# dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X847 dvss.t219 a_4921_n3946# a_5346_n3990# dvss.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X848 a_n12731_9395# a_n13109_1995# avss.t303 sky130_fd_pr__res_xhigh_po_1p41 l=35
X849 comparator_0.vt vin.t106 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X850 schmitt_trigger_0.in.t9 dvss.t117 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X851 rstring_mux_0.vtrip6.t0 rstring_mux_0.otrip_decoded_avdd[6] vin.t17 avss.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X852 avdd.t386 rstring_mux_0.ena_b rstring_mux_0.vtop.t1 avdd.t385 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X853 dvdd.t113 a_10874_n1026# a_10874_n2222# dvdd.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X854 avdd.t94 avdd.t93 avdd.t94 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=8
X855 dvss.t500 schmitt_trigger_0.out.t13 sky130_fd_sc_hd__inv_4_0.Y dvss.t499 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X856 dvss.t254 a_429_n1142# a_1636_n1478# dvss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X857 avdd.t7 a_n5907_n2876# a_n5214_n3990# avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X858 a_n22549_n11914# a_n22927_n15834# avss.t275 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X859 vin.t31 avdd.t91 vin.t31 avdd.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X860 rstring_mux_0.otrip_decoded_avdd[4] a_n2588_n3212# dvss.t543 dvss.t542 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X861 rstring_mux_0.otrip_decoded_b_avdd[8] rstring_mux_0.otrip_decoded_avdd[8] avdd.t198 avdd.t197 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X862 rstring_mux_0.otrip_decoded_b_avdd[3] rstring_mux_0.otrip_decoded_avdd[3] avdd.t37 avdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X863 a_5346_n3990# a_4921_n3946# dvss.t217 dvss.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X864 schmitt_trigger_0.m.t6 schmitt_trigger_0.in.t10 dvdd.t23 dvdd.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X865 dvdd.t25 schmitt_trigger_0.in.t11 schmitt_trigger_0.m.t7 dvdd.t24 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X866 ibias_gen_0.vn1.t8 ibias_gen_0.isrc_sel_b avss.t359 avss.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X867 avss.t89 avss.t88 avss.t89 avss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X868 dvss.t311 a_10515_n1026# a_10874_n1026# dvss.t310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X869 avdd.t333 ibias_gen_0.ena rstring_mux_0.ena_b avdd.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X870 vin.t68 avss.t86 vin.t68 avss.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X871 a_n7429_n11914# a_n7807_n15834# avss.t297 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X872 dvss.t126 a_7033_n3946# a_7458_n3990# dvss.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X873 comparator_0.vnn vbg_1v2.t23 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X874 rstring_mux_0.otrip_decoded_avdd[1] a_n6812_n1478# dvss.t110 dvss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X875 vin.t30 avdd.t89 vin.t30 avdd.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X876 a_n8195_9395# a_n8573_1995# avss.t335 sky130_fd_pr__res_xhigh_po_1p41 l=35
X877 ovout.t0 sky130_fd_sc_hd__inv_4_0.Y dvss.t148 dvss.t147 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X878 vin.t67 avss.t84 vin.t67 avss.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X879 rstring_mux_0.otrip_decoded_b_avdd[12] rstring_mux_0.otrip_decoded_avdd[12] avdd.t271 avdd.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X880 comparator_0.vn comparator_0.ena_b avss.t180 avss.t179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X881 comparator_0.vpp vin.t107 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X882 rstring_mux_0.otrip_decoded_avdd[7] a_n476_n1478# avdd.t285 avdd.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X883 vin.t66 avss.t82 vin.t66 avss.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X884 avdd.t314 a_n8019_n2876# a_n7326_n3990# avdd.t313 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X885 comparator_0.vt avss.t398 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X886 a_2809_n3946# a_2441_n2964# dvss.t333 dvss.t332 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X887 a_5423_n11914# a_5801_n15834# avss.t382 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X888 vin.t65 avss.t80 vin.t65 avss.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X889 dvss.t443 a_n3527_n3946# a_n3102_n3990# dvss.t442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X890 ibg_200n ibias_gen_0.ena_b a_n15529_n2223# avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X891 schmitt_trigger_0.out.t3 schmitt_trigger_0.m.t17 dvss.t381 dvss.t380 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X892 dvss.t37 a_9145_n3946# a_9570_n3990# dvss.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X893 rstring_mux_0.vtrip1.t5 rstring_mux_0.vtrip2.t5 avss.t383 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X894 avdd.t219 comparator_0.vnn comparator_0.vpp avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X895 avdd.t88 avdd.t86 avdd.t87 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=8
X896 avdd.t85 avdd.t83 avdd.t85 avdd.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=8
X897 a_n26329_n11914# a_n26707_n15834# avss.t280 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X898 a_n3102_n3990# a_n3527_n3946# dvss.t441 dvss.t440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X899 rstring_mux_0.vtrip11.t4 rstring_mux_0.otrip_decoded_avdd[11] vin.t81 avss.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X900 dvss.t1 a_n3795_n2876# a_n2588_n3212# dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X901 a_7033_n3946# a_6665_n2964# dvss.t417 dvss.t416 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X902 ovout.t16 sky130_fd_sc_hd__inv_4_0.Y dvdd.t29 dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X903 schmitt_trigger_0.in.t12 dvss.t118 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X904 dvss.t525 a_n5639_n3946# a_n5214_n3990# dvss.t524 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X905 comparator_0.vnn comparator_0.vpp avdd.t15 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X906 rstring_mux_0.vtrip14.t2 rstring_mux_0.otrip_decoded_avdd[14] vin.t24 avss.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X907 dvss.t401 a_4553_n2964# a_4653_n2876# dvss.t400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X908 avss.t247 comparator_0.vm comparator_0.vm avss.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X909 dvss.t379 otrip_decoded[6].t1 a_n1783_n2964# dvss.t378 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X910 rstring_mux_0.vtrip11.t0 rstring_mux_0.vtrip10.t2 avss.t22 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X911 comparator_0.vpp vin.t108 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X912 rstring_mux_0.vtrip9.t3 rstring_mux_0.otrip_decoded_b_avdd[9] vin.t49 avdd.t309 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X913 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t14 dvdd.t63 dvdd.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X914 avss.t79 avss.t77 avss.t79 avss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X915 comparator_0.vt avss.t399 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X916 a_n21793_n11914# a_n21415_n15834# avss.t263 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X917 schmitt_trigger_0.in.t13 dvss.t119 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X918 a_n5214_n3990# a_n5639_n3946# dvss.t523 dvss.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X919 avdd.t372 a_n1683_n1142# a_n476_n1478# avdd.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X920 rstring_mux_0.otrip_decoded_b_avdd[10] rstring_mux_0.otrip_decoded_avdd[10] avss.t12 avss.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X921 comparator_0.vt vbg_1v2.t24 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X922 dvss.t3 a_n5907_n2876# a_n4700_n3212# dvss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X923 vin.t4 rstring_mux_0.otrip_decoded_b_avdd[3] rstring_mux_0.vtrip3.t3 avdd.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X924 dcomp comparator_0.n1 avss.t29 avss.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X925 a_n5917_n11914# a_n6295_n15834# avss.t258 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X926 a_9145_n3946# a_8777_n2964# dvss.t321 dvss.t320 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X927 a_1122_n3990# a_697_n3946# dvss.t284 dvss.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X928 avdd.t331 a_n990_n2256# a_n1683_n1142# avdd.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X929 vin.t64 avss.t75 vin.t64 avss.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X930 dvss.t478 a_n7751_n3946# a_n7326_n3990# dvss.t477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X931 ibias_gen_0.vn0.t18 ibias_gen_0.vp0.t13 avdd.t369 avdd.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X932 avss.t74 avss.t71 avss.t73 avss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X933 comparator_0.vt vin.t109 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X934 schmitt_trigger_0.in.t14 dvss.t120 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X935 dvss.t377 otrip_decoded[4].t1 a_n3895_n2964# dvss.t376 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X936 avdd.t82 avdd.t79 avdd.t81 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X937 ibias_gen_0.vr.t2 avss.t69 ibias_gen_0.ve.t4 avss.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X938 vin.t63 avss.t67 vin.t63 avss.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X939 a_697_n3946# a_329_n2964# dvss.t184 dvss.t183 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X940 avdd.t53 comparator_0.n1 dcomp avdd.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X941 ibias_gen_0.vp0.t7 avss.t65 ibias_gen_0.vn0.t5 avss.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X942 rstring_mux_0.otrip_decoded_avdd[12] a_5860_n3212# dvss.t122 dvss.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X943 ibias_gen_0.vn1.t1 avdd.t77 ibias_gen_0.vp1.t0 avdd.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X944 avdd.t13 comparator_0.vpp comparator_0.vnn avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X945 vin.t93 avss.t63 vin.t93 avss.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X946 avss.t27 comparator_0.n1 dcomp avss.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X947 avss.t62 avss.t60 avss.t62 avss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X948 dvss.t365 a_n8019_n2876# a_n6812_n3212# dvss.t364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X949 avdd.t1 a_n3795_n2876# a_n3102_n3990# avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X950 comparator_0.vnn comparator_0.vnn avdd.t218 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X951 a_429_n2876# a_329_n2964# dvss.t182 dvss.t181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X952 a_3234_n3990# a_2809_n3946# dvss.t196 dvss.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X953 schmitt_trigger_0.m.t9 schmitt_trigger_0.out.t15 dvdd.t61 dvdd.t60 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X954 comparator_0.vt avss.t400 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X955 a_n24817_n11914# a_n25195_n15834# avss.t334 sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X956 a_10874_n1026# a_10874_n2222# dvdd.t132 dvdd.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
X957 rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.otrip_decoded_avdd[6] avss.t195 avss.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X958 dvss.t383 otrip_decoded[2].t1 a_n6007_n2964# dvss.t382 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X959 ibias_gen_0.vstart.t1 vbg_1v2.t25 ibias_gen_0.vn0.t16 avss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X960 dvss.t215 a_4921_n3946# a_5346_n3990# dvss.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X961 dvss.t85 a_429_n2876# a_1636_n3212# dvss.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
R0 vin.n80 vin.n79 63.7962
R1 vin.n20 vin.t20 53.91
R2 vin.n128 vin.t92 51.0275
R3 vin.n136 vin.n2 48.371
R4 vin.n6 vin.n5 48.371
R5 vin.n23 vin.n22 48.371
R6 vin.n27 vin.n26 48.371
R7 vin.n31 vin.n30 48.371
R8 vin.n35 vin.n34 48.371
R9 vin.n39 vin.n38 48.371
R10 vin.n43 vin.n42 48.371
R11 vin.n47 vin.n46 48.371
R12 vin.n51 vin.n50 48.371
R13 vin.n55 vin.n54 48.371
R14 vin.n59 vin.n58 48.371
R15 vin.n63 vin.n62 48.371
R16 vin.n83 vin.n82 48.371
R17 vin.n133 vin.n0 48.371
R18 vin.n135 vin.n134 45.4885
R19 vin.n4 vin.n3 45.4885
R20 vin.n8 vin.n7 45.4885
R21 vin.n21 vin.n9 45.4885
R22 vin.n25 vin.n10 45.4885
R23 vin.n29 vin.n11 45.4885
R24 vin.n33 vin.n12 45.4885
R25 vin.n37 vin.n13 45.4885
R26 vin.n41 vin.n14 45.4885
R27 vin.n45 vin.n15 45.4885
R28 vin.n49 vin.n16 45.4885
R29 vin.n53 vin.n17 45.4885
R30 vin.n57 vin.n18 45.4885
R31 vin.n61 vin.n19 45.4885
R32 vin.n85 vin.n84 45.4885
R33 vin.n86 vin.t69 21.0726
R34 vin.n129 vin.t10 20.2802
R35 vin.n132 vin.n127 17.7666
R36 vin.n125 vin.n124 17.7666
R37 vin.n122 vin.n121 17.7666
R38 vin.n119 vin.n118 17.7666
R39 vin.n116 vin.n115 17.7666
R40 vin.n113 vin.n112 17.7666
R41 vin.n110 vin.n109 17.7666
R42 vin.n107 vin.n106 17.7666
R43 vin.n104 vin.n103 17.7666
R44 vin.n101 vin.n100 17.7666
R45 vin.n98 vin.n97 17.7666
R46 vin.n95 vin.n94 17.7666
R47 vin.n92 vin.n91 17.7666
R48 vin.n89 vin.n88 17.7666
R49 vin.n130 vin.n129 17.7666
R50 vin.n132 vin.n131 16.9742
R51 vin.n126 vin.n125 16.9742
R52 vin.n123 vin.n122 16.9742
R53 vin.n120 vin.n119 16.9742
R54 vin.n117 vin.n116 16.9742
R55 vin.n114 vin.n113 16.9742
R56 vin.n111 vin.n110 16.9742
R57 vin.n108 vin.n107 16.9742
R58 vin.n105 vin.n104 16.9742
R59 vin.n102 vin.n101 16.9742
R60 vin.n99 vin.n98 16.9742
R61 vin.n96 vin.n95 16.9742
R62 vin.n93 vin.n92 16.9742
R63 vin.n90 vin.n89 16.9742
R64 vin.n87 vin.n86 16.9742
R65 vin.n78 vin.t94 13.1361
R66 vin.n76 vin.t95 13.1361
R67 vin.n74 vin.t106 13.1361
R68 vin.n72 vin.t109 13.1361
R69 vin.n70 vin.t105 13.1361
R70 vin.n68 vin.t102 13.1361
R71 vin.n66 vin.t103 13.1361
R72 vin.n65 vin.t101 13.1361
R73 vin.n78 vin.t99 11.2285
R74 vin.n76 vin.t100 11.2285
R75 vin.n74 vin.t97 11.2285
R76 vin.n72 vin.t98 11.2285
R77 vin.n70 vin.t96 11.2285
R78 vin.n68 vin.t107 11.2285
R79 vin.n66 vin.t108 11.2285
R80 vin.n65 vin.t104 11.2285
R81 vin.n134 vin.t78 5.5395
R82 vin.n134 vin.t84 5.5395
R83 vin.n2 vin.t83 5.5395
R84 vin.t30 vin.n2 5.5395
R85 vin.n3 vin.t30 5.5395
R86 vin.n3 vin.t7 5.5395
R87 vin.n6 vin.t6 5.5395
R88 vin.t71 vin.n6 5.5395
R89 vin.n7 vin.t71 5.5395
R90 vin.n7 vin.t15 5.5395
R91 vin.n22 vin.t14 5.5395
R92 vin.n22 vin.t76 5.5395
R93 vin.t76 vin.n21 5.5395
R94 vin.n21 vin.t52 5.5395
R95 vin.n26 vin.t51 5.5395
R96 vin.n26 vin.t74 5.5395
R97 vin.t74 vin.n25 5.5395
R98 vin.n25 vin.t56 5.5395
R99 vin.n30 vin.t55 5.5395
R100 vin.n30 vin.t32 5.5395
R101 vin.t32 vin.n29 5.5395
R102 vin.n29 vin.t50 5.5395
R103 vin.n34 vin.t49 5.5395
R104 vin.n34 vin.t41 5.5395
R105 vin.t41 vin.n33 5.5395
R106 vin.n33 vin.t57 5.5395
R107 vin.n38 vin.t58 5.5395
R108 vin.n38 vin.t39 5.5395
R109 vin.t39 vin.n37 5.5395
R110 vin.n37 vin.t59 5.5395
R111 vin.n42 vin.t60 5.5395
R112 vin.n42 vin.t73 5.5395
R113 vin.t73 vin.n41 5.5395
R114 vin.n41 vin.t86 5.5395
R115 vin.n46 vin.t85 5.5395
R116 vin.n46 vin.t75 5.5395
R117 vin.t75 vin.n45 5.5395
R118 vin.n45 vin.t53 5.5395
R119 vin.n50 vin.t54 5.5395
R120 vin.n50 vin.t77 5.5395
R121 vin.t77 vin.n49 5.5395
R122 vin.n49 vin.t89 5.5395
R123 vin.n54 vin.t90 5.5395
R124 vin.n54 vin.t40 5.5395
R125 vin.t40 vin.n53 5.5395
R126 vin.n53 vin.t4 5.5395
R127 vin.n58 vin.t5 5.5395
R128 vin.n58 vin.t42 5.5395
R129 vin.t42 vin.n57 5.5395
R130 vin.n57 vin.t61 5.5395
R131 vin.n62 vin.t62 5.5395
R132 vin.n62 vin.t72 5.5395
R133 vin.t72 vin.n61 5.5395
R134 vin.n61 vin.t48 5.5395
R135 vin.n83 vin.t47 5.5395
R136 vin.t31 vin.n83 5.5395
R137 vin.n84 vin.t31 5.5395
R138 vin.n84 vin.t21 5.5395
R139 vin.n133 vin.t91 5.5395
R140 vin.t78 vin.n133 5.5395
R141 vin.n67 vin.n65 5.04858
R142 vin.n67 vin.n66 4.5005
R143 vin.n69 vin.n68 4.5005
R144 vin.n71 vin.n70 4.5005
R145 vin.n73 vin.n72 4.5005
R146 vin.n75 vin.n74 4.5005
R147 vin.n77 vin.n76 4.5005
R148 vin.n79 vin.n78 4.5005
R149 vin vin.n0 3.76065
R150 vin.n80 vin.n20 3.4105
R151 vin.n82 vin.n81 3.4105
R152 vin.n64 vin.n63 3.4105
R153 vin.n60 vin.n59 3.4105
R154 vin.n56 vin.n55 3.4105
R155 vin.n52 vin.n51 3.4105
R156 vin.n48 vin.n47 3.4105
R157 vin.n44 vin.n43 3.4105
R158 vin.n40 vin.n39 3.4105
R159 vin.n36 vin.n35 3.4105
R160 vin.n32 vin.n31 3.4105
R161 vin.n28 vin.n27 3.4105
R162 vin.n24 vin.n23 3.4105
R163 vin.n5 vin.n1 3.4105
R164 vin.n137 vin.n136 3.4105
R165 vin.n131 vin.t64 3.3065
R166 vin.n131 vin.t25 3.3065
R167 vin.n127 vin.t24 3.3065
R168 vin.n127 vin.t44 3.3065
R169 vin.t44 vin.n126 3.3065
R170 vin.n126 vin.t80 3.3065
R171 vin.n124 vin.t79 3.3065
R172 vin.n124 vin.t46 3.3065
R173 vin.t46 vin.n123 3.3065
R174 vin.n123 vin.t26 3.3065
R175 vin.n121 vin.t27 3.3065
R176 vin.n121 vin.t36 3.3065
R177 vin.t36 vin.n120 3.3065
R178 vin.n120 vin.t82 3.3065
R179 vin.n118 vin.t81 3.3065
R180 vin.n118 vin.t45 3.3065
R181 vin.t45 vin.n117 3.3065
R182 vin.n117 vin.t2 3.3065
R183 vin.n115 vin.t3 3.3065
R184 vin.n115 vin.t43 3.3065
R185 vin.t43 vin.n114 3.3065
R186 vin.n114 vin.t22 3.3065
R187 vin.n112 vin.t23 3.3065
R188 vin.n112 vin.t33 3.3065
R189 vin.t33 vin.n111 3.3065
R190 vin.n111 vin.t13 3.3065
R191 vin.n109 vin.t12 3.3065
R192 vin.n109 vin.t67 3.3065
R193 vin.t67 vin.n108 3.3065
R194 vin.n108 vin.t38 3.3065
R195 vin.n106 vin.t37 3.3065
R196 vin.n106 vin.t93 3.3065
R197 vin.t93 vin.n105 3.3065
R198 vin.n105 vin.t16 3.3065
R199 vin.n103 vin.t17 3.3065
R200 vin.n103 vin.t65 3.3065
R201 vin.t65 vin.n102 3.3065
R202 vin.n102 vin.t18 3.3065
R203 vin.n100 vin.t19 3.3065
R204 vin.n100 vin.t68 3.3065
R205 vin.t68 vin.n99 3.3065
R206 vin.n99 vin.t9 3.3065
R207 vin.n97 vin.t8 3.3065
R208 vin.n97 vin.t63 3.3065
R209 vin.t63 vin.n96 3.3065
R210 vin.n96 vin.t0 3.3065
R211 vin.n94 vin.t1 3.3065
R212 vin.n94 vin.t35 3.3065
R213 vin.t35 vin.n93 3.3065
R214 vin.n93 vin.t29 3.3065
R215 vin.n91 vin.t28 3.3065
R216 vin.n91 vin.t66 3.3065
R217 vin.t66 vin.n90 3.3065
R218 vin.n90 vin.t88 3.3065
R219 vin.n88 vin.t87 3.3065
R220 vin.n88 vin.t34 3.3065
R221 vin.t34 vin.n87 3.3065
R222 vin.n87 vin.t70 3.3065
R223 vin.n130 vin.t11 3.3065
R224 vin.t64 vin.n130 3.3065
R225 vin.n135 vin.n132 1.98319
R226 vin.n125 vin.n4 1.98319
R227 vin.n122 vin.n8 1.98319
R228 vin.n119 vin.n9 1.98319
R229 vin.n116 vin.n10 1.98319
R230 vin.n113 vin.n11 1.98319
R231 vin.n110 vin.n12 1.98319
R232 vin.n107 vin.n13 1.98319
R233 vin.n104 vin.n14 1.98319
R234 vin.n101 vin.n15 1.98319
R235 vin.n98 vin.n16 1.98319
R236 vin.n95 vin.n17 1.98319
R237 vin.n92 vin.n18 1.98319
R238 vin.n89 vin.n19 1.98319
R239 vin.n86 vin.n85 1.98319
R240 vin.n129 vin.n128 1.98319
R241 vin.n69 vin.n67 0.548577
R242 vin.n71 vin.n69 0.548577
R243 vin.n73 vin.n71 0.548577
R244 vin.n75 vin.n73 0.548577
R245 vin.n77 vin.n75 0.548577
R246 vin.n79 vin.n77 0.548577
R247 vin.n81 vin.n80 0.384333
R248 vin.n81 vin.n64 0.384333
R249 vin.n64 vin.n60 0.384333
R250 vin.n60 vin.n56 0.384333
R251 vin.n56 vin.n52 0.384333
R252 vin.n52 vin.n48 0.384333
R253 vin.n48 vin.n44 0.384333
R254 vin.n44 vin.n40 0.384333
R255 vin.n40 vin.n36 0.384333
R256 vin.n36 vin.n32 0.384333
R257 vin.n32 vin.n28 0.384333
R258 vin.n28 vin.n24 0.384333
R259 vin.n24 vin.n1 0.384333
R260 vin.n137 vin.n1 0.384333
R261 vin vin.n137 0.0341833
R262 vin.n136 vin.n135 0.00218919
R263 vin.n5 vin.n4 0.00218919
R264 vin.n23 vin.n8 0.00218919
R265 vin.n27 vin.n9 0.00218919
R266 vin.n31 vin.n10 0.00218919
R267 vin.n35 vin.n11 0.00218919
R268 vin.n39 vin.n12 0.00218919
R269 vin.n43 vin.n13 0.00218919
R270 vin.n47 vin.n14 0.00218919
R271 vin.n51 vin.n15 0.00218919
R272 vin.n55 vin.n16 0.00218919
R273 vin.n59 vin.n17 0.00218919
R274 vin.n63 vin.n18 0.00218919
R275 vin.n82 vin.n19 0.00218919
R276 vin.n85 vin.n20 0.00218919
R277 vin.n128 vin.n0 0.00218919
R278 rstring_mux_0.vtrip12.n2 rstring_mux_0.vtrip12.n0 50.7022
R279 rstring_mux_0.vtrip12.n3 rstring_mux_0.vtrip12.n2 18.1477
R280 rstring_mux_0.vtrip12.n2 rstring_mux_0.vtrip12.n1 13.8791
R281 rstring_mux_0.vtrip12.n3 rstring_mux_0.vtrip12.t5 10.6297
R282 rstring_mux_0.vtrip12.n0 rstring_mux_0.vtrip12.t1 5.5395
R283 rstring_mux_0.vtrip12.n0 rstring_mux_0.vtrip12.t0 5.5395
R284 rstring_mux_0.vtrip12.n1 rstring_mux_0.vtrip12.t3 3.3065
R285 rstring_mux_0.vtrip12.n1 rstring_mux_0.vtrip12.t4 3.3065
R286 rstring_mux_0.vtrip12.t2 rstring_mux_0.vtrip12.n3 0.826075
R287 avss.n761 avss.n14 128525
R288 avss.n14 avss.n12 128525
R289 avss.n13 avss.n12 128525
R290 avss.n761 avss.n13 128525
R291 avss.n662 avss.n355 98666.5
R292 avss.n655 avss.n355 70225
R293 avss.n267 avss.n26 68021.9
R294 avss.n332 avss.n326 45524.4
R295 avss.n332 avss.n327 45524.4
R296 avss.n677 avss.n327 45524.4
R297 avss.n677 avss.n326 45524.4
R298 avss.n435 avss.n390 45524.4
R299 avss.n439 avss.n390 45524.4
R300 avss.n435 avss.n391 45524.4
R301 avss.n439 avss.n391 45524.4
R302 avss.n149 avss.n26 45183
R303 avss.n436 avss.n427 35028.6
R304 avss.n729 avss.n309 21059.4
R305 avss.n731 avss.n309 21059.4
R306 avss.n731 avss.n308 21059.4
R307 avss.n729 avss.n308 21059.4
R308 avss.t211 avss.n355 20202
R309 avss.n449 avss.n360 18174.6
R310 avss.n651 avss.n360 18174.6
R311 avss.n449 avss.n361 18174.6
R312 avss.n651 avss.n361 18174.6
R313 avss.n747 avss.n24 16300.9
R314 avss.n744 avss.n24 16300.9
R315 avss.n747 avss.n25 16300.9
R316 avss.n744 avss.n25 16300.9
R317 avss.n267 avss.n266 12588.9
R318 avss.n664 avss.n341 12517.1
R319 avss.n664 avss.n342 12517.1
R320 avss.n350 avss.n342 12517.1
R321 avss.n350 avss.n341 12517.1
R322 avss.n662 avss.n661 10118.5
R323 avss.n760 avss.n15 8350.87
R324 avss.n755 avss.n16 8350.87
R325 avss.n755 avss.n15 8350.87
R326 avss.n759 avss.n16 8341.08
R327 avss.n518 avss.n514 7742.83
R328 avss.n520 avss.n514 7742.83
R329 avss.n519 avss.n518 7742.83
R330 avss.n520 avss.n519 7742.83
R331 avss.n683 avss.n325 7610.36
R332 avss.n684 avss.n325 7610.36
R333 avss.n684 avss.n324 7610.36
R334 avss.n683 avss.n324 7610.36
R335 avss.n663 avss.n662 6546.95
R336 avss.n407 avss.n396 5644.38
R337 avss.n407 avss.n397 5644.38
R338 avss.n418 avss.n397 5644.38
R339 avss.n418 avss.n396 5644.38
R340 avss.n517 avss.n512 4175.68
R341 avss.n521 avss.n512 4175.68
R342 avss.n517 avss.n513 4175.68
R343 avss.n521 avss.n513 4175.68
R344 avss.n446 avss.n384 4139.43
R345 avss.n453 avss.n384 4139.43
R346 avss.n453 avss.n385 4139.43
R347 avss.n446 avss.n385 4139.43
R348 avss.n656 avss.n357 3978.07
R349 avss.n660 avss.n357 3978.07
R350 avss.n660 avss.n356 3978.07
R351 avss.n656 avss.n356 3978.07
R352 avss.t78 avss.t186 3966.94
R353 avss.t186 avss.t192 3966.94
R354 avss.t190 avss.t188 3966.94
R355 avss.t188 avss.t96 3966.94
R356 avss.n421 avss.n392 3902.33
R357 avss.n421 avss.n393 3902.33
R358 avss.n425 avss.n393 3902.33
R359 avss.n425 avss.n392 3902.33
R360 avss.n268 avss.n3 2998.14
R361 avss.n674 avss.n673 2957.93
R362 avss.n434 avss.n433 2957.93
R363 avss.n434 avss.n429 2940.24
R364 avss.n673 avss.n331 2935.34
R365 avss.n260 avss.n259 2905.02
R366 avss.n45 avss.n44 2905.02
R367 avss.n246 avss.n245 2905.02
R368 avss.n61 avss.n60 2905.02
R369 avss.n232 avss.n231 2905.02
R370 avss.n77 avss.n76 2905.02
R371 avss.n218 avss.n217 2905.02
R372 avss.n93 avss.n92 2905.02
R373 avss.n204 avss.n203 2905.02
R374 avss.n109 avss.n108 2905.02
R375 avss.n190 avss.n189 2905.02
R376 avss.n125 avss.n124 2905.02
R377 avss.n176 avss.n175 2905.02
R378 avss.n141 avss.n140 2905.02
R379 avss.n162 avss.n161 2905.02
R380 avss.n763 avss.n762 2538.7
R381 avss.t26 avss.n384 2436.62
R382 avss.t211 avss.n385 2436.62
R383 avss.n732 avss.n307 2366.87
R384 avss.n732 avss.n306 2366.87
R385 avss.n433 avss.n389 2361.98
R386 avss.n728 avss.n306 2344.28
R387 avss.n728 avss.n307 2344.28
R388 avss.n450 avss.t78 2304.08
R389 avss.n652 avss.t96 2304.08
R390 avss.n564 avss.n548 2087.09
R391 avss.n589 avss.n538 2084.98
R392 avss.n648 avss.n364 2054.02
R393 avss.n640 avss.n364 2054.02
R394 avss.n428 avss.n388 2048.38
R395 avss.n582 avss.n580 2039.85
R396 avss.n606 avss.n605 2039.84
R397 avss.t192 avss.n448 1983.47
R398 avss.n448 avss.t190 1983.47
R399 avss.t44 avss.t120 1910.53
R400 avss.t45 avss.t44 1910.53
R401 avss.t43 avss.t25 1910.53
R402 avss.t91 avss.t43 1910.53
R403 avss.n640 avss.n363 1894.78
R404 avss.n649 avss.n648 1894.78
R405 avss.n743 avss.n269 1813.84
R406 avss.n765 avss.n10 1735.47
R407 avss.n766 avss.n10 1735.47
R408 avss.n766 avss.n9 1735.47
R409 avss.n765 avss.n9 1735.47
R410 avss.n353 avss.t45 1647.77
R411 avss.n749 avss.n22 1602.64
R412 avss.n676 avss.n328 1487.81
R413 avss.n676 avss.n675 1487.81
R414 avss.n331 avss.n328 1439.24
R415 avss.n675 avss.n674 1439.24
R416 avss.n665 avss.n340 1435.48
R417 avss.n349 avss.n340 1435.48
R418 avss.n775 avss.n3 1414.29
R419 avss.n666 avss.n339 1385.79
R420 avss.n348 avss.n339 1385.79
R421 avss.n447 avss.t30 1301
R422 avss.t34 avss.n447 1301
R423 avss.t120 avss.n350 1286.14
R424 avss.n663 avss.t91 1253.64
R425 avss.t34 avss.t36 1081.77
R426 avss.t28 avss.t26 1081.77
R427 avss.t32 avss.t28 1081.77
R428 avss.t38 avss.t32 1081.77
R429 avss.t30 avss.t38 1081.77
R430 avss.t36 avss.t40 1081.77
R431 avss.t40 avss.t209 1081.77
R432 avss.t25 avss.n354 1008.7
R433 avss.n516 avss.n509 976.942
R434 avss.n516 avss.n515 976.942
R435 avss.n523 avss.n522 976.188
R436 avss.n522 avss.n511 974.683
R437 avss.n26 avss.n3 939.895
R438 avss.n452 avss.t30 925.769
R439 avss.n452 avss.t34 925.769
R440 avss.n354 avss.t70 901.822
R441 avss.n451 avss.t211 887.293
R442 avss.n682 avss.n681 874.542
R443 avss.n682 avss.n322 874.542
R444 avss.n260 avss.n30 815.444
R445 avss.n44 avss.n41 815.444
R446 avss.n247 avss.n246 815.444
R447 avss.n60 avss.n57 815.444
R448 avss.n233 avss.n232 815.444
R449 avss.n76 avss.n73 815.444
R450 avss.n219 avss.n218 815.444
R451 avss.n92 avss.n89 815.444
R452 avss.n205 avss.n204 815.444
R453 avss.n108 avss.n105 815.444
R454 avss.n191 avss.n190 815.444
R455 avss.n124 avss.n121 815.444
R456 avss.n177 avss.n176 815.444
R457 avss.n140 avss.n137 815.444
R458 avss.n163 avss.n162 815.444
R459 avss.n149 avss.n148 815.444
R460 avss.n273 avss.n23 796.612
R461 avss.n273 avss.n272 782.683
R462 avss.n777 avss.n776 769.572
R463 avss.n686 avss.n685 765.741
R464 avss.n685 avss.n323 765.741
R465 avss.n742 avss.n270 759.718
R466 avss.n266 avss.t150 755.986
R467 avss.n259 avss.t228 755.986
R468 avss.t362 avss.n45 755.986
R469 avss.n245 avss.t233 755.986
R470 avss.t367 avss.n61 755.986
R471 avss.n231 avss.t11 755.986
R472 avss.t222 avss.n77 755.986
R473 avss.n217 avss.t157 755.986
R474 avss.t267 avss.n93 755.986
R475 avss.n203 avss.t194 755.986
R476 avss.t201 avss.n109 755.986
R477 avss.n189 avss.t51 755.986
R478 avss.t8 avss.n125 755.986
R479 avss.n175 avss.t240 755.986
R480 avss.t373 avss.n141 755.986
R481 avss.n161 avss.t347 755.986
R482 avss.t323 avss.t321 731.963
R483 avss.t179 avss.t183 731.963
R484 avss.t183 avss.n653 684.673
R485 avss.t321 avss.n654 668.225
R486 avss.n417 avss.n398 649.788
R487 avss.n408 avss.n398 649.788
R488 avss.n581 avss.t114 625.516
R489 avss.n588 avss.t114 625.516
R490 avss.t114 avss.n532 614.321
R491 avss.n599 avss.t114 614.321
R492 avss.n655 avss.t323 602.431
R493 avss.n271 avss.n270 598.966
R494 avss.t114 avss.n571 598.606
R495 avss.n572 avss.t114 598.606
R496 avss.n440 avss.n389 595.953
R497 avss.n557 avss.t114 588.343
R498 avss.n555 avss.t114 588.343
R499 avss.n578 avss.n577 585
R500 avss.n576 avss.n545 585
R501 avss.n545 avss.n544 585
R502 avss.n575 avss.n574 585
R503 avss.n574 avss.n573 585
R504 avss.n547 avss.n546 585
R505 avss.n572 avss.n547 585
R506 avss.n570 avss.n569 585
R507 avss.n571 avss.n570 585
R508 avss.n568 avss.n549 585
R509 avss.n549 avss.n548 585
R510 avss.n567 avss.n566 585
R511 avss.n551 avss.n550 585
R512 avss.n593 avss.n592 585
R513 avss.n590 avss.n540 585
R514 avss.n590 avss.n589 585
R515 avss.n587 avss.n586 585
R516 avss.n588 avss.n587 585
R517 avss.n585 avss.n541 585
R518 avss.n581 avss.n541 585
R519 avss.n584 avss.n583 585
R520 avss.n583 avss.n582 585
R521 avss.n543 avss.n542 585
R522 avss.n594 avss.n539 585
R523 avss.n596 avss.n595 585
R524 avss.n597 avss.n596 585
R525 avss.n537 avss.n536 585
R526 avss.n598 avss.n537 585
R527 avss.n601 avss.n600 585
R528 avss.n600 avss.n599 585
R529 avss.n602 avss.n534 585
R530 avss.n534 avss.n532 585
R531 avss.n604 avss.n603 585
R532 avss.n605 avss.n604 585
R533 avss.n535 avss.n533 585
R534 avss.n529 avss.n527 585
R535 avss.n562 avss.n561 585
R536 avss.n563 avss.n562 585
R537 avss.n560 avss.n553 585
R538 avss.n553 avss.n552 585
R539 avss.n559 avss.n558 585
R540 avss.n558 avss.n557 585
R541 avss.n556 avss.n554 585
R542 avss.n556 avss.n555 585
R543 avss.n528 avss.n526 585
R544 avss.n530 avss.n528 585
R545 avss.n609 avss.n608 585
R546 avss.n608 avss.n607 585
R547 avss.n774 avss.n773 585
R548 avss.n775 avss.n774 585
R549 avss.n2 avss.n1 585
R550 avss.n265 avss.n264 585
R551 avss.n266 avss.n265 585
R552 avss.n263 avss.n27 585
R553 avss.n30 avss.n27 585
R554 avss.n262 avss.n261 585
R555 avss.n261 avss.n260 585
R556 avss.n258 avss.n257 585
R557 avss.n259 avss.n258 585
R558 avss.n32 avss.n31 585
R559 avss.n41 avss.n31 585
R560 avss.n43 avss.n42 585
R561 avss.n44 avss.n43 585
R562 avss.n250 avss.n38 585
R563 avss.n45 avss.n38 585
R564 avss.n249 avss.n248 585
R565 avss.n248 avss.n247 585
R566 avss.n40 avss.n39 585
R567 avss.n246 avss.n40 585
R568 avss.n244 avss.n243 585
R569 avss.n245 avss.n244 585
R570 avss.n47 avss.n46 585
R571 avss.n57 avss.n46 585
R572 avss.n59 avss.n58 585
R573 avss.n60 avss.n59 585
R574 avss.n236 avss.n54 585
R575 avss.n61 avss.n54 585
R576 avss.n235 avss.n234 585
R577 avss.n234 avss.n233 585
R578 avss.n56 avss.n55 585
R579 avss.n232 avss.n56 585
R580 avss.n230 avss.n229 585
R581 avss.n231 avss.n230 585
R582 avss.n63 avss.n62 585
R583 avss.n73 avss.n62 585
R584 avss.n75 avss.n74 585
R585 avss.n76 avss.n75 585
R586 avss.n222 avss.n70 585
R587 avss.n77 avss.n70 585
R588 avss.n221 avss.n220 585
R589 avss.n220 avss.n219 585
R590 avss.n72 avss.n71 585
R591 avss.n218 avss.n72 585
R592 avss.n216 avss.n215 585
R593 avss.n217 avss.n216 585
R594 avss.n79 avss.n78 585
R595 avss.n89 avss.n78 585
R596 avss.n91 avss.n90 585
R597 avss.n92 avss.n91 585
R598 avss.n208 avss.n86 585
R599 avss.n93 avss.n86 585
R600 avss.n207 avss.n206 585
R601 avss.n206 avss.n205 585
R602 avss.n88 avss.n87 585
R603 avss.n204 avss.n88 585
R604 avss.n202 avss.n201 585
R605 avss.n203 avss.n202 585
R606 avss.n95 avss.n94 585
R607 avss.n105 avss.n94 585
R608 avss.n107 avss.n106 585
R609 avss.n108 avss.n107 585
R610 avss.n194 avss.n102 585
R611 avss.n109 avss.n102 585
R612 avss.n193 avss.n192 585
R613 avss.n192 avss.n191 585
R614 avss.n104 avss.n103 585
R615 avss.n190 avss.n104 585
R616 avss.n188 avss.n187 585
R617 avss.n189 avss.n188 585
R618 avss.n111 avss.n110 585
R619 avss.n121 avss.n110 585
R620 avss.n123 avss.n122 585
R621 avss.n124 avss.n123 585
R622 avss.n180 avss.n118 585
R623 avss.n125 avss.n118 585
R624 avss.n179 avss.n178 585
R625 avss.n178 avss.n177 585
R626 avss.n120 avss.n119 585
R627 avss.n176 avss.n120 585
R628 avss.n174 avss.n173 585
R629 avss.n175 avss.n174 585
R630 avss.n127 avss.n126 585
R631 avss.n137 avss.n126 585
R632 avss.n139 avss.n138 585
R633 avss.n140 avss.n139 585
R634 avss.n166 avss.n134 585
R635 avss.n141 avss.n134 585
R636 avss.n165 avss.n164 585
R637 avss.n164 avss.n163 585
R638 avss.n136 avss.n135 585
R639 avss.n162 avss.n136 585
R640 avss.n160 avss.n159 585
R641 avss.n161 avss.n160 585
R642 avss.n143 avss.n142 585
R643 avss.n148 avss.n142 585
R644 avss.n151 avss.n150 585
R645 avss.n150 avss.n149 585
R646 avss.n441 avss.n388 584.659
R647 avss.n409 avss.n399 540.989
R648 avss.n416 avss.n399 540.989
R649 avss.n160 avss.n142 539.294
R650 avss.n150 avss.n142 539.294
R651 avss.n164 avss.n134 539.294
R652 avss.n164 avss.n136 539.294
R653 avss.n174 avss.n126 539.294
R654 avss.n139 avss.n126 539.294
R655 avss.n178 avss.n118 539.294
R656 avss.n178 avss.n120 539.294
R657 avss.n188 avss.n110 539.294
R658 avss.n123 avss.n110 539.294
R659 avss.n192 avss.n102 539.294
R660 avss.n192 avss.n104 539.294
R661 avss.n202 avss.n94 539.294
R662 avss.n107 avss.n94 539.294
R663 avss.n206 avss.n86 539.294
R664 avss.n206 avss.n88 539.294
R665 avss.n216 avss.n78 539.294
R666 avss.n91 avss.n78 539.294
R667 avss.n220 avss.n70 539.294
R668 avss.n220 avss.n72 539.294
R669 avss.n230 avss.n62 539.294
R670 avss.n75 avss.n62 539.294
R671 avss.n234 avss.n54 539.294
R672 avss.n234 avss.n56 539.294
R673 avss.n244 avss.n46 539.294
R674 avss.n59 avss.n46 539.294
R675 avss.n248 avss.n38 539.294
R676 avss.n248 avss.n40 539.294
R677 avss.n258 avss.n31 539.294
R678 avss.n43 avss.n31 539.294
R679 avss.n265 avss.n27 539.294
R680 avss.n261 avss.n27 539.294
R681 avss.n774 avss.n2 539.294
R682 avss.n3 avss.t326 492.382
R683 avss.n454 avss.n383 477.741
R684 avss.n445 avss.n383 477.741
R685 avss.n661 avss.t181 474.954
R686 avss.n657 avss.n359 459.295
R687 avss.n658 avss.n657 459.295
R688 avss.n659 avss.n658 459.295
R689 avss.n558 avss.n556 456.416
R690 avss.n600 avss.n534 456.416
R691 avss.n587 avss.n541 456.416
R692 avss.n570 avss.n547 456.416
R693 avss.n424 avss.n394 425.264
R694 avss.n422 avss.n394 420.43
R695 avss.n423 avss.n422 420.43
R696 avss.n424 avss.n423 420.43
R697 avss.n444 avss.n382 401.812
R698 avss.n455 avss.n382 401.812
R699 avss.n321 avss.t65 392.769
R700 avss.n401 avss.t133 392.692
R701 avss.n402 avss.t106 392.664
R702 avss.n21 avss.t75 384.515
R703 avss.n277 avss.t129 384.515
R704 avss.n279 avss.t122 384.515
R705 avss.n280 avss.t131 384.515
R706 avss.n281 avss.t127 384.515
R707 avss.n282 avss.t104 384.515
R708 avss.n283 avss.t84 384.515
R709 avss.n285 avss.t63 384.515
R710 avss.n287 avss.t86 384.515
R711 avss.n288 avss.t67 384.515
R712 avss.n289 avss.t115 384.515
R713 avss.n290 avss.t82 384.515
R714 avss.n291 avss.t108 384.515
R715 avss.n278 avss.t135 384.454
R716 avss.n286 avss.t80 384.454
R717 avss.n582 avss.n581 363.548
R718 avss.n589 avss.n588 363.548
R719 avss.n605 avss.n532 357.041
R720 avss.n599 avss.n598 357.041
R721 avss.n598 avss.n597 357.041
R722 avss.n597 avss.n538 357.041
R723 avss.n571 avss.n548 347.908
R724 avss.n573 avss.n572 347.908
R725 avss.n573 avss.n544 347.908
R726 avss.n580 avss.n544 347.908
R727 avss.n564 avss.n563 341.943
R728 avss.n563 avss.n552 341.943
R729 avss.n557 avss.n552 341.943
R730 avss.n555 avss.n530 341.943
R731 avss.n607 avss.n530 341.943
R732 avss.n607 avss.n606 341.943
R733 avss.n451 avss.n450 340.805
R734 avss.n494 avss.n481 333.334
R735 avss.n489 avss.n488 333.334
R736 avss.n504 avss.n479 333.334
R737 avss.t342 avss.n11 323.332
R738 avss.t342 avss.n763 323.332
R739 avss.n362 avss.n358 318.495
R740 avss.n441 avss.n440 302.307
R741 avss.n11 avss.n3 301.202
R742 avss.t19 avss.t56 298.923
R743 avss.t56 avss.t258 298.923
R744 avss.t258 avss.t331 298.923
R745 avss.t331 avss.t55 298.923
R746 avss.t55 avss.t152 298.923
R747 avss.t152 avss.t297 298.923
R748 avss.t297 avss.t328 298.923
R749 avss.t328 avss.t312 298.923
R750 avss.n591 avss.n538 283.521
R751 avss.n580 avss.n579 283.521
R752 avss.n743 avss.n742 274.072
R753 avss.n748 avss.n23 270.683
R754 avss.t70 avss.n353 262.753
R755 avss.n565 avss.n564 262.719
R756 avss.n606 avss.n531 262.719
R757 avss.n749 avss.n748 238.306
R758 avss.n653 avss.n652 227.298
R759 avss.n745 avss.t298 211.297
R760 avss.t137 avss.n394 209.756
R761 avss.n423 avss.t137 209.756
R762 avss.n272 avss.n271 208.189
R763 avss.n764 avss.n8 202.918
R764 avss.n767 avss.n8 202.918
R765 avss.n776 avss.n775 200.215
R766 avss.n268 avss.t19 199.304
R767 avss.t209 avss.n451 194.476
R768 avss.n764 avss.n7 193.918
R769 avss.n768 avss.n767 186.73
R770 avss.n499 avss.n498 185
R771 avss.n500 avss.n486 185
R772 avss.n492 avss.n491 185
R773 avss.n493 avss.n481 185
R774 avss.t113 avss.n481 185
R775 avss.n495 avss.n494 185
R776 avss.n497 avss.n496 185
R777 avss.n488 avss.n487 185
R778 avss.n490 avss.n489 185
R779 avss.n480 avss.n478 185
R780 avss.n505 avss.n504 185
R781 avss.n504 avss.t113 185
R782 avss.n479 avss.n477 185
R783 avss.n502 avss.n501 185
R784 avss.n776 avss.n2 184.572
R785 avss.t335 avss.t274 170.34
R786 avss.t361 avss.t335 170.34
R787 avss.t153 avss.t361 170.34
R788 avss.t304 avss.t153 170.34
R789 avss.t330 avss.t304 170.34
R790 avss.t21 avss.t330 170.34
R791 avss.t332 avss.t42 170.34
R792 avss.t214 avss.t332 170.34
R793 avss.t46 avss.t345 170.34
R794 avss.t254 avss.t46 170.34
R795 avss.t303 avss.t254 170.34
R796 avss.t251 avss.t303 170.34
R797 avss.t281 avss.t251 170.34
R798 avss.t272 avss.t281 170.34
R799 avss.t207 avss.t272 170.34
R800 avss.t220 avss.t207 170.34
R801 avss.t6 avss.t220 170.34
R802 avss.n438 avss.n355 166.736
R803 avss.n650 avss.n363 159.248
R804 avss.n650 avss.n649 159.248
R805 avss.t48 avss.t317 155.921
R806 avss.t378 avss.t317 155.921
R807 avss.t357 avss.t378 155.921
R808 avss.t58 avss.t357 155.921
R809 avss.t23 avss.t58 155.921
R810 avss.t300 avss.t277 155.921
R811 avss.t154 avss.t300 155.921
R812 avss.t337 avss.t154 155.921
R813 avss.t376 avss.t337 155.921
R814 avss.t306 avss.t376 155.921
R815 avss.t237 avss.t306 155.921
R816 avss.t296 avss.t237 155.921
R817 avss.t271 avss.t296 155.921
R818 avss.t242 avss.t271 155.921
R819 avss.t262 avss.t242 155.921
R820 avss.t261 avss.t262 155.921
R821 avss.t270 avss.t261 155.921
R822 avss.t216 avss.t270 155.921
R823 avss.t382 avss.t216 155.921
R824 avss.t257 avss.t382 155.921
R825 avss.t354 avss.t257 155.921
R826 avss.t318 avss.t354 155.921
R827 avss.t4 avss.t318 155.921
R828 avss.n155 avss.t348 149.067
R829 avss.n146 avss.t374 149.067
R830 avss.n169 avss.t241 149.067
R831 avss.n130 avss.t9 149.067
R832 avss.n183 avss.t52 149.067
R833 avss.n114 avss.t202 149.067
R834 avss.n197 avss.t195 149.067
R835 avss.n98 avss.t268 149.067
R836 avss.n211 avss.t158 149.067
R837 avss.n82 avss.t223 149.067
R838 avss.n225 avss.t12 149.067
R839 avss.n66 avss.t368 149.067
R840 avss.n239 avss.t234 149.067
R841 avss.n50 avss.t363 149.067
R842 avss.n253 avss.t229 149.067
R843 avss.n34 avss.t151 149.067
R844 avss.n4 avss.t327 149.067
R845 avss.t336 avss.t23 142.516
R846 avss.n746 avss.t148 140.655
R847 avss.n562 avss.n553 132.635
R848 avss.n558 avss.n553 132.635
R849 avss.n556 avss.n528 132.635
R850 avss.n608 avss.n528 132.635
R851 avss.n604 avss.n533 132.635
R852 avss.n604 avss.n534 132.635
R853 avss.n600 avss.n537 132.635
R854 avss.n596 avss.n537 132.635
R855 avss.n596 avss.n539 132.635
R856 avss.n583 avss.n543 132.635
R857 avss.n583 avss.n541 132.635
R858 avss.n590 avss.n587 132.635
R859 avss.n592 avss.n590 132.635
R860 avss.n566 avss.n549 132.635
R861 avss.n570 avss.n549 132.635
R862 avss.n574 avss.n547 132.635
R863 avss.n574 avss.n545 132.635
R864 avss.n578 avss.n545 132.635
R865 avss.t311 avss.t185 120.487
R866 avss.t208 avss.t282 120.487
R867 avss.t341 avss.t230 120.487
R868 avss.t230 avss.t20 120.487
R869 avss.t274 avss.n435 119.504
R870 avss.n762 avss.t312 117.829
R871 avss.n384 avss.n382 117.001
R872 avss.n385 avss.n383 117.001
R873 avss.n657 avss.n656 117.001
R874 avss.n656 avss.n655 117.001
R875 avss.n660 avss.n659 117.001
R876 avss.n661 avss.n660 117.001
R877 avss.n765 avss.n764 117.001
R878 avss.t342 avss.n765 117.001
R879 avss.n767 avss.n766 117.001
R880 avss.n766 avss.t342 117.001
R881 avss.n438 avss.t6 114.462
R882 avss.t277 avss.n13 113.772
R883 avss.n436 avss.t21 113.561
R884 avss.t349 avss.t244 113.532
R885 avss.t2 avss.t310 113.475
R886 avss.n491 avss.n481 113.334
R887 avss.n504 avss.n480 113.334
R888 avss.t149 avss.t76 112.272
R889 avss.t227 avss.t226 112.272
R890 avss.t130 avss.t365 112.272
R891 avss.t364 avss.t136 112.272
R892 avss.t232 avss.t235 112.272
R893 avss.t123 avss.t369 112.272
R894 avss.t369 avss.t366 112.272
R895 avss.t132 avss.t13 112.272
R896 avss.t14 avss.t128 112.272
R897 avss.t221 avss.t224 112.272
R898 avss.t105 avss.t155 112.272
R899 avss.t156 avss.t85 112.272
R900 avss.t266 avss.t269 112.272
R901 avss.t64 avss.t197 112.272
R902 avss.t196 avss.t81 112.272
R903 avss.t81 avss.t200 112.272
R904 avss.t203 avss.t87 112.272
R905 avss.t50 avss.t49 112.272
R906 avss.t68 avss.t7 112.272
R907 avss.t10 avss.t116 112.272
R908 avss.t239 avss.t238 112.272
R909 avss.t83 avss.t372 112.272
R910 avss.t371 avss.t109 112.272
R911 avss.t350 avss.t349 112.272
R912 avss.t340 avss.t203 109.749
R913 avss.t264 avss.t132 108.487
R914 avss.n427 avss.t336 105.188
R915 avss.t235 avss.t53 102.18
R916 avss.t259 avss.t0 101.999
R917 avss.t197 avss.t351 100.918
R918 avss.t109 avss.t276 99.6565
R919 avss.n659 avss.n358 99.0123
R920 avss.n9 avss.n7 97.5005
R921 avss.n11 avss.n9 97.5005
R922 avss.n10 avss.n8 97.5005
R923 avss.n763 avss.n10 97.5005
R924 avss.t16 avss.t50 95.8721
R925 avss.t217 avss.t14 94.6106
R926 avss.n762 avss.t48 94.46
R927 avss.t20 avss.n14 89.9625
R928 avss.t136 avss.t165 88.3032
R929 avss.n373 avss.t27 88.2028
R930 avss.n377 avss.t212 88.2028
R931 avss.n613 avss.t182 88.2028
R932 avss.t161 avss.t198 87.975
R933 avss.n615 avss.t322 87.8727
R934 avss.n486 avss.n484 87.6787
R935 avss.n498 avss.n484 87.6787
R936 avss.n614 avss.t180 87.5075
R937 avss.n613 avss.t184 87.5075
R938 avss.t269 avss.t255 87.0418
R939 avss.n681 avss.n323 86.2123
R940 avss.n686 avss.n322 86.2123
R941 avss.n417 avss.n416 86.2123
R942 avss.n409 avss.n408 86.2123
R943 avss.t372 avss.t260 85.7803
R944 avss.n437 avss.t214 85.1705
R945 avss.t345 avss.n437 85.1705
R946 avss.n769 avss.t343 85.1191
R947 avss.n631 avss.t126 82.9912
R948 avss.n629 avss.t98 82.9912
R949 avss.n463 avss.t100 82.9912
R950 avss.t79 avss.n458 82.9912
R951 avss.n363 avss.n362 82.824
R952 avss.n649 avss.n358 82.824
R953 avss.t375 avss.t68 81.9959
R954 avss.t380 avss.t218 81.2813
R955 avss.t314 avss.t17 81.2813
R956 avss.t308 avss.t206 81.2813
R957 avss.t263 avss.t339 81.2813
R958 avss.t377 avss.t253 81.2813
R959 avss.t24 avss.t204 81.2813
R960 avss.t275 avss.t315 81.2813
R961 avss.t338 avss.t199 81.2813
R962 avss.t381 avss.t219 81.2813
R963 avss.t177 avss.t178 81.2813
R964 avss.t252 avss.t334 81.2813
R965 avss.t352 avss.t47 81.2813
R966 avss.t305 avss.t370 81.2813
R967 avss.t319 avss.t245 81.2813
R968 avss.t15 avss.t280 81.2813
R969 avss.t59 avss.t205 81.2813
R970 avss.t309 avss.t273 81.2813
R971 avss.t355 avss.n351 80.9625
R972 avss.t22 avss.t221 80.7344
R973 avss.t333 avss.t149 79.473
R974 avss.t282 avss.n678 78.7313
R975 avss.t113 avss.n482 77.7851
R976 avss.t113 avss.n483 77.7851
R977 avss.t346 avss.t358 76.5001
R978 avss.n420 avss.t61 76.1813
R979 avss.n426 avss.t316 75.2251
R980 avss.t365 avss.t256 74.4271
R981 avss.t85 avss.t279 73.1656
R982 avss.t238 avss.t302 71.9042
R983 avss.n375 avss.n374 70.9775
R984 avss.n373 avss.n372 70.9775
R985 avss.n379 avss.n378 70.9775
R986 avss.n377 avss.n376 70.9775
R987 avss.n638 avss.n637 70.9612
R988 avss.n636 avss.n635 70.9612
R989 avss.n644 avss.n643 70.9612
R990 avss.n646 avss.n645 70.9612
R991 avss.n462 avss.n461 70.9612
R992 avss.n460 avss.n459 70.9612
R993 avss.t113 avss.n485 70.8113
R994 avss.t113 avss.n503 70.8113
R995 avss.n498 avss.n497 70.0005
R996 avss.n502 avss.n486 70.0005
R997 avss.t383 avss.t10 68.1198
R998 avss.t379 avss.t324 67.8939
R999 avss.n353 avss.t54 67.2564
R1000 avss.t384 avss.t105 66.8583
R1001 avss.n404 avss.t57 65.9814
R1002 avss.t265 avss.t227 65.5968
R1003 avss.t138 avss.n395 64.7064
R1004 avss.n679 avss.t208 63.7501
R1005 avss.n654 avss.t179 63.7388
R1006 avss.n680 avss.t236 62.4751
R1007 avss.t226 avss.t344 60.551
R1008 avss.t307 avss.n352 60.2439
R1009 avss.n746 avss.n267 59.9202
R1010 avss.n533 avss.n531 59.5655
R1011 avss.n566 avss.n565 59.5655
R1012 avss.n565 avss.n551 59.5655
R1013 avss.n531 avss.n529 59.5655
R1014 avss.n30 avss.t150 59.46
R1015 avss.n41 avss.t228 59.46
R1016 avss.n247 avss.t362 59.46
R1017 avss.n57 avss.t233 59.46
R1018 avss.n233 avss.t367 59.46
R1019 avss.n73 avss.t11 59.46
R1020 avss.n219 avss.t222 59.46
R1021 avss.n89 avss.t157 59.46
R1022 avss.n205 avss.t267 59.46
R1023 avss.n105 avss.t194 59.46
R1024 avss.n191 avss.t201 59.46
R1025 avss.n121 avss.t51 59.46
R1026 avss.n177 avss.t8 59.46
R1027 avss.n137 avss.t240 59.46
R1028 avss.n163 avss.t373 59.46
R1029 avss.n148 avss.t347 59.46
R1030 avss.t155 avss.t246 59.2895
R1031 avss.t116 avss.t313 58.028
R1032 avss.t147 avss.n680 58.0127
R1033 avss.n343 avss.t69 57.0602
R1034 avss.t42 avss.n436 56.7805
R1035 avss.t163 avss.t320 56.7377
R1036 avss.t164 avss.t107 56.7377
R1037 avss.t174 avss.t66 56.7377
R1038 avss.t173 avss.t171 56.7377
R1039 avss.t170 avss.t168 56.7377
R1040 avss.t167 avss.t166 56.7377
R1041 avss.t169 avss.t172 56.7377
R1042 avss.t236 avss.n679 56.7377
R1043 avss.t168 avss.t225 55.7814
R1044 avss.t231 avss.n404 54.5064
R1045 avss.t313 avss.t239 54.2436
R1046 avss.t166 avss.t72 53.5502
R1047 avss.n406 avss.n405 53.2314
R1048 avss.n651 avss.n650 53.1823
R1049 avss.n652 avss.n651 53.1823
R1050 avss.n449 avss.n364 53.1823
R1051 avss.n450 avss.n449 53.1823
R1052 avss.t246 avss.t156 52.9822
R1053 avss.t324 avss.t353 52.594
R1054 avss.t344 avss.t130 51.7207
R1055 avss.t176 avss.t169 50.6815
R1056 avss.n445 avss.n444 49.8123
R1057 avss.n455 avss.n454 49.8123
R1058 avss.n757 avss.n756 49.4893
R1059 avss.n758 avss.n757 49.4335
R1060 avss.t171 avss.t215 48.769
R1061 avss.t113 avss.n484 48.6621
R1062 avss.n653 avss.t181 47.2902
R1063 avss.t76 avss.t265 46.6748
R1064 avss.n756 avss.n754 45.4402
R1065 avss.t224 avss.t384 45.4133
R1066 avss.t185 avss.n426 45.2627
R1067 avss.n394 avss.n392 45.0005
R1068 avss.t138 avss.n392 45.0005
R1069 avss.n423 avss.n393 45.0005
R1070 avss.t138 avss.n393 45.0005
R1071 avss.t7 avss.t383 44.1519
R1072 avss.n494 avss.n485 43.3803
R1073 avss.n503 avss.n479 43.3803
R1074 avss.n497 avss.n485 43.3803
R1075 avss.n503 avss.n502 43.3803
R1076 avss.t18 avss.t174 41.7565
R1077 avss.n678 avss.t243 41.7565
R1078 avss.n730 avss.t213 41.4378
R1079 avss.t302 avss.t83 40.3675
R1080 avss.n18 avss.n17 40.092
R1081 avss.n406 avss.t346 39.2065
R1082 avss.t218 avss.t243 39.2065
R1083 avss.t17 avss.t380 39.2065
R1084 avss.t206 avss.t314 39.2065
R1085 avss.t339 avss.t308 39.2065
R1086 avss.t253 avss.t263 39.2065
R1087 avss.t204 avss.t377 39.2065
R1088 avss.t315 avss.t24 39.2065
R1089 avss.t199 avss.t275 39.2065
R1090 avss.t329 avss.t338 39.2065
R1091 avss.t54 avss.t307 39.2065
R1092 avss.t301 avss.t381 39.2065
R1093 avss.t219 avss.t177 39.2065
R1094 avss.t178 avss.t252 39.2065
R1095 avss.t334 avss.t352 39.2065
R1096 avss.t47 avss.t305 39.2065
R1097 avss.t370 avss.t319 39.2065
R1098 avss.t245 avss.t15 39.2065
R1099 avss.t280 avss.t59 39.2065
R1100 avss.t205 avss.t309 39.2065
R1101 avss.t273 avss.t355 39.2065
R1102 avss.t279 avss.t266 39.106
R1103 avss.t256 avss.t364 37.8445
R1104 avss.n159 avss.n143 36.1417
R1105 avss.n151 avss.n143 36.1417
R1106 avss.n166 avss.n165 36.1417
R1107 avss.n165 avss.n135 36.1417
R1108 avss.n173 avss.n127 36.1417
R1109 avss.n138 avss.n127 36.1417
R1110 avss.n180 avss.n179 36.1417
R1111 avss.n179 avss.n119 36.1417
R1112 avss.n187 avss.n111 36.1417
R1113 avss.n122 avss.n111 36.1417
R1114 avss.n194 avss.n193 36.1417
R1115 avss.n193 avss.n103 36.1417
R1116 avss.n201 avss.n95 36.1417
R1117 avss.n106 avss.n95 36.1417
R1118 avss.n208 avss.n207 36.1417
R1119 avss.n207 avss.n87 36.1417
R1120 avss.n215 avss.n79 36.1417
R1121 avss.n90 avss.n79 36.1417
R1122 avss.n222 avss.n221 36.1417
R1123 avss.n221 avss.n71 36.1417
R1124 avss.n229 avss.n63 36.1417
R1125 avss.n74 avss.n63 36.1417
R1126 avss.n236 avss.n235 36.1417
R1127 avss.n235 avss.n55 36.1417
R1128 avss.n243 avss.n47 36.1417
R1129 avss.n58 avss.n47 36.1417
R1130 avss.n250 avss.n249 36.1417
R1131 avss.n249 avss.n39 36.1417
R1132 avss.n257 avss.n32 36.1417
R1133 avss.n42 avss.n32 36.1417
R1134 avss.n264 avss.n263 36.1417
R1135 avss.n263 avss.n262 36.1417
R1136 avss.n773 avss.n1 36.1417
R1137 avss.n777 avss.n1 36.1417
R1138 avss.n269 avss.n22 36.1417
R1139 avss.t107 avss.t295 36.019
R1140 avss.t285 avss.t134 35.7003
R1141 avss.n495 avss.n493 35.5561
R1142 avss.n490 avss.n487 35.5561
R1143 avss.n562 avss.n551 35.1094
R1144 avss.n608 avss.n529 35.1094
R1145 avss.t5 avss.t360 34.744
R1146 avss.n744 avss.n743 34.4123
R1147 avss.n745 avss.n744 34.4123
R1148 avss.n748 avss.n747 34.4123
R1149 avss.n747 avss.n746 34.4123
R1150 avss.t148 avss.t333 32.7987
R1151 avss.t310 avss.t161 32.5128
R1152 avss.n350 avss.n349 32.5005
R1153 avss.n665 avss.n664 32.5005
R1154 avss.n664 avss.n663 32.5005
R1155 avss.n425 avss.n424 32.5005
R1156 avss.n426 avss.n425 32.5005
R1157 avss.n422 avss.n421 32.5005
R1158 avss.n421 avss.n420 32.5005
R1159 avss.n418 avss.n417 32.5005
R1160 avss.n419 avss.n418 32.5005
R1161 avss.n408 avss.n407 32.5005
R1162 avss.n407 avss.n406 32.5005
R1163 avss.n681 avss.n324 32.5005
R1164 avss.n405 avss.n324 32.5005
R1165 avss.n325 avss.n322 32.5005
R1166 avss.n680 avss.n325 32.5005
R1167 avss.t128 avss.t22 31.5372
R1168 avss.t49 avss.t375 30.2757
R1169 avss.n569 avss.n546 29.6559
R1170 avss.n586 avss.n585 29.6559
R1171 avss.n602 avss.n601 29.6559
R1172 avss.t353 avss.t138 29.6441
R1173 avss.n491 avss.n482 29.4328
R1174 avss.n488 avss.n483 29.4328
R1175 avss.n489 avss.n482 29.4328
R1176 avss.n483 avss.n480 29.4328
R1177 avss.t134 avss.t299 29.0066
R1178 avss.n362 avss.n359 28.9887
R1179 avss.n405 avss.t213 28.0503
R1180 avss.n419 avss.t198 27.7316
R1181 avss.t299 avss.t164 27.7316
R1182 avss.t244 avss.n745 27.1221
R1183 avss.n666 avss.n665 27.1064
R1184 avss.n349 avss.n348 27.1064
R1185 avss.n617 avss.n612 26.6319
R1186 avss.t260 avss.t371 26.4913
R1187 avss.n296 avss.t110 26.4633
R1188 avss.n303 avss.t88 26.4633
R1189 avss.n691 avss.t101 26.4633
R1190 avss.n697 avss.t117 26.4633
R1191 avss.n704 avss.t142 26.4633
R1192 avss.n710 avss.t60 26.4633
R1193 avss.n720 avss.t139 26.4633
R1194 avss.n715 avss.t145 26.4633
R1195 avss.n318 avss.t71 26.4633
R1196 avss.n313 avss.t93 26.4633
R1197 avss.t358 avss.t283 25.8191
R1198 avss.t255 avss.t64 25.2299
R1199 avss.n335 avss.t90 25.2191
R1200 avss.n344 avss.t119 25.2191
R1201 avss.t165 avss.t232 23.9684
R1202 avss.n400 avss.t160 23.7186
R1203 avss.n411 avss.t359 23.4728
R1204 avss.n414 avss.t162 23.4728
R1205 avss.n400 avss.t325 23.4728
R1206 avss.n359 avss.n356 22.5005
R1207 avss.n654 avss.n356 22.5005
R1208 avss.n658 avss.n357 22.5005
R1209 avss.n654 avss.n357 22.5005
R1210 avss.t66 avss.t5 21.9941
R1211 avss.n432 avss.n431 21.1018
R1212 avss.t360 avss.t285 21.0379
R1213 avss.n352 avss.t301 21.0379
R1214 avss.n431 avss.n430 20.9741
R1215 avss.n446 avss.n445 20.8934
R1216 avss.n447 avss.n446 20.8934
R1217 avss.n454 avss.n453 20.8934
R1218 avss.n453 avss.n452 20.8934
R1219 avss.t295 avss.t163 20.7191
R1220 avss.n300 avss.n299 20.3733
R1221 avss.n302 avss.n301 20.3733
R1222 avss.n694 avss.n693 20.3733
R1223 avss.n696 avss.n695 20.3733
R1224 avss.n707 avss.n706 20.3733
R1225 avss.n709 avss.n708 20.3733
R1226 avss.n719 avss.n718 20.3733
R1227 avss.n717 avss.n716 20.3733
R1228 avss.n317 avss.n316 20.3733
R1229 avss.n315 avss.n314 20.3733
R1230 avss avss.n499 20.2672
R1231 avss.n398 avss.n396 20.1729
R1232 avss.n404 avss.n396 20.1729
R1233 avss.n399 avss.n397 20.1729
R1234 avss.n404 avss.n397 20.1729
R1235 avss.n413 avss.n412 20.1668
R1236 avss.t0 avss.t231 18.4879
R1237 avss.t283 avss.t259 18.1691
R1238 avss.n296 avss.t112 18.0193
R1239 avss.n303 avss.t89 18.0193
R1240 avss.n691 avss.t103 18.0193
R1241 avss.n697 avss.t118 18.0193
R1242 avss.n704 avss.t144 18.0193
R1243 avss.n710 avss.t62 18.0193
R1244 avss.n720 avss.t141 18.0193
R1245 avss.t146 avss.n715 18.0193
R1246 avss.n318 avss.t74 18.0193
R1247 avss.t94 avss.n313 18.0193
R1248 avss.n592 avss.n591 17.9618
R1249 avss.n579 avss.n543 17.9618
R1250 avss.n579 avss.n578 17.9618
R1251 avss.n591 avss.n539 17.9618
R1252 avss.n506 avss.n505 17.9561
R1253 avss.n429 avss.n428 17.6946
R1254 avss.t13 avss.t217 17.6611
R1255 avss.n506 avss.n477 17.6005
R1256 avss.n395 avss.t159 17.5317
R1257 avss.n335 avss.t92 17.2863
R1258 avss.n344 avss.t121 17.2863
R1259 avss.n432 avss.n387 17.0331
R1260 avss.n559 avss 16.7292
R1261 avss.n374 avss.t39 16.5305
R1262 avss.n374 avss.t31 16.5305
R1263 avss.n372 avss.t29 16.5305
R1264 avss.n372 avss.t33 16.5305
R1265 avss.n378 avss.t35 16.5305
R1266 avss.n378 avss.t37 16.5305
R1267 avss.n376 avss.t41 16.5305
R1268 avss.n376 avss.t210 16.5305
R1269 avss.n637 avss.t250 16.5305
R1270 avss.n637 avss.t125 16.5305
R1271 avss.n635 avss.t189 16.5305
R1272 avss.n635 avss.t97 16.5305
R1273 avss.n643 avss.t248 16.5305
R1274 avss.n643 avss.t247 16.5305
R1275 avss.n645 avss.t193 16.5305
R1276 avss.n645 avss.t191 16.5305
R1277 avss.t100 avss.n462 16.5305
R1278 avss.n462 avss.t249 16.5305
R1279 avss.n459 avss.t79 16.5305
R1280 avss.n459 avss.t187 16.5305
R1281 avss.t87 avss.t16 16.3996
R1282 avss.n469 avss.t399 15.9785
R1283 avss.n470 avss.t400 15.9785
R1284 avss.n471 avss.t397 15.9785
R1285 avss.n472 avss.t398 15.9785
R1286 avss.n473 avss.t396 15.9785
R1287 avss.n474 avss.t391 15.9785
R1288 avss.n475 avss.t392 15.9785
R1289 avss.n476 avss.t388 15.9785
R1290 avss.n420 avss.t379 15.9379
R1291 avss.n627 avss.t394 15.8834
R1292 avss.n626 avss.t395 15.8834
R1293 avss.n625 avss.t390 15.8834
R1294 avss.n624 avss.t393 15.8834
R1295 avss.n623 avss.t389 15.8834
R1296 avss.n622 avss.t386 15.8834
R1297 avss.n621 avss.t387 15.8834
R1298 avss.n620 avss.t385 15.8834
R1299 avss.n427 avss.t311 15.3004
R1300 avss.n500 avss 15.2894
R1301 avss.t173 avss.t18 14.9817
R1302 avss.n403 avss.n323 14.9605
R1303 avss.n416 avss.n415 14.9605
R1304 avss.n410 avss.n409 14.9605
R1305 avss.n687 avss.n686 14.9605
R1306 avss.n430 avss.n386 14.8972
R1307 avss.n753 avss.n752 14.0996
R1308 avss.n631 avss.t124 14.0925
R1309 avss.n629 avss.t95 14.0925
R1310 avss.n463 avss.t99 14.0925
R1311 avss.n458 avss.t77 14.0925
R1312 avss.n353 avss.t329 14.0254
R1313 avss.t172 avss.t147 13.0692
R1314 avss.n554 avss 12.9272
R1315 avss.n683 avss.n682 12.7179
R1316 avss.t173 avss.n683 12.7179
R1317 avss.n685 avss.n684 12.7179
R1318 avss.n684 avss.t173 12.7179
R1319 avss.t276 avss.t350 12.6152
R1320 avss.n671 avss.n293 12.189
R1321 avss.n496 avss.n495 12.0894
R1322 avss.n493 avss.n492 12.0894
R1323 avss.n501 avss.n477 12.0894
R1324 avss.n505 avss.n478 12.0894
R1325 avss.n669 avss.t356 11.9874
R1326 avss.n753 avss.t278 11.9517
R1327 avss.n769 avss.n768 11.8447
R1328 avss.t351 avss.t196 11.3537
R1329 avss.n444 avss.n443 10.3105
R1330 avss.n456 avss.n455 10.3105
R1331 avss.t53 avss.t123 10.0922
R1332 avss.n760 avss.n759 9.78874
R1333 avss.n628 avss.n627 9.59836
R1334 avss.n469 avss.n468 9.57265
R1335 avss.n758 avss.n17 9.42238
R1336 avss.n734 avss.n733 9.42076
R1337 avss.n733 avss.n305 9.42076
R1338 avss.n275 avss.n271 9.35869
R1339 avss.n274 avss.n273 9.35222
R1340 avss.n23 avss.n19 9.34791
R1341 avss.n276 avss.n270 9.33929
R1342 avss.n742 avss.n741 9.33929
R1343 avss.n772 avss.n4 9.30641
R1344 avss.n35 avss.n34 9.3005
R1345 avss.n34 avss.n33 9.3005
R1346 avss.n253 avss.n252 9.3005
R1347 avss.n254 avss.n253 9.3005
R1348 avss.n51 avss.n50 9.3005
R1349 avss.n50 avss.n49 9.3005
R1350 avss.n239 avss.n238 9.3005
R1351 avss.n240 avss.n239 9.3005
R1352 avss.n67 avss.n66 9.3005
R1353 avss.n66 avss.n65 9.3005
R1354 avss.n225 avss.n224 9.3005
R1355 avss.n226 avss.n225 9.3005
R1356 avss.n83 avss.n82 9.3005
R1357 avss.n82 avss.n81 9.3005
R1358 avss.n211 avss.n210 9.3005
R1359 avss.n212 avss.n211 9.3005
R1360 avss.n99 avss.n98 9.3005
R1361 avss.n98 avss.n97 9.3005
R1362 avss.n197 avss.n196 9.3005
R1363 avss.n198 avss.n197 9.3005
R1364 avss.n115 avss.n114 9.3005
R1365 avss.n114 avss.n113 9.3005
R1366 avss.n183 avss.n182 9.3005
R1367 avss.n184 avss.n183 9.3005
R1368 avss.n131 avss.n130 9.3005
R1369 avss.n130 avss.n129 9.3005
R1370 avss.n169 avss.n168 9.3005
R1371 avss.n170 avss.n169 9.3005
R1372 avss.n147 avss.n146 9.3005
R1373 avss.n146 avss.n145 9.3005
R1374 avss.n155 avss.n154 9.3005
R1375 avss.n156 avss.n155 9.3005
R1376 avss.n257 avss.n256 9.3005
R1377 avss.n255 avss.n32 9.3005
R1378 avss.n42 avss.n36 9.3005
R1379 avss.n251 avss.n250 9.3005
R1380 avss.n249 avss.n37 9.3005
R1381 avss.n48 avss.n39 9.3005
R1382 avss.n243 avss.n242 9.3005
R1383 avss.n241 avss.n47 9.3005
R1384 avss.n58 avss.n52 9.3005
R1385 avss.n237 avss.n236 9.3005
R1386 avss.n235 avss.n53 9.3005
R1387 avss.n64 avss.n55 9.3005
R1388 avss.n229 avss.n228 9.3005
R1389 avss.n227 avss.n63 9.3005
R1390 avss.n74 avss.n68 9.3005
R1391 avss.n223 avss.n222 9.3005
R1392 avss.n221 avss.n69 9.3005
R1393 avss.n80 avss.n71 9.3005
R1394 avss.n215 avss.n214 9.3005
R1395 avss.n213 avss.n79 9.3005
R1396 avss.n90 avss.n84 9.3005
R1397 avss.n209 avss.n208 9.3005
R1398 avss.n207 avss.n85 9.3005
R1399 avss.n96 avss.n87 9.3005
R1400 avss.n201 avss.n200 9.3005
R1401 avss.n199 avss.n95 9.3005
R1402 avss.n106 avss.n100 9.3005
R1403 avss.n195 avss.n194 9.3005
R1404 avss.n193 avss.n101 9.3005
R1405 avss.n112 avss.n103 9.3005
R1406 avss.n187 avss.n186 9.3005
R1407 avss.n185 avss.n111 9.3005
R1408 avss.n122 avss.n116 9.3005
R1409 avss.n181 avss.n180 9.3005
R1410 avss.n179 avss.n117 9.3005
R1411 avss.n128 avss.n119 9.3005
R1412 avss.n173 avss.n172 9.3005
R1413 avss.n171 avss.n127 9.3005
R1414 avss.n138 avss.n132 9.3005
R1415 avss.n167 avss.n166 9.3005
R1416 avss.n165 avss.n133 9.3005
R1417 avss.n144 avss.n135 9.3005
R1418 avss.n159 avss.n158 9.3005
R1419 avss.n157 avss.n143 9.3005
R1420 avss.n152 avss.n151 9.3005
R1421 avss.n264 avss.n20 9.3005
R1422 avss.n263 avss.n28 9.3005
R1423 avss.n262 avss.n29 9.3005
R1424 avss.n667 avss.n666 9.3005
R1425 avss.n348 avss.n347 9.3005
R1426 avss.n333 avss.n328 9.3005
R1427 avss.n675 avss.n294 9.3005
R1428 avss.n442 avss.n441 9.3005
R1429 avss.n5 avss.n4 9.3005
R1430 avss.n773 avss.n772 9.3005
R1431 avss.n1 avss.n0 9.3005
R1432 avss.n778 avss.n777 9.3005
R1433 avss.n750 avss.n749 9.3005
R1434 avss.n739 avss.n738 9.20927
R1435 avss.n16 avss.n14 9.0005
R1436 avss.n15 avss.n13 9.0005
R1437 avss.n672 avss.n670 8.81442
R1438 avss.n567 avss.n550 8.61832
R1439 avss.n568 avss.n567 8.61832
R1440 avss.n569 avss.n568 8.61832
R1441 avss.n575 avss.n546 8.61832
R1442 avss.n576 avss.n575 8.61832
R1443 avss.n577 avss.n576 8.61832
R1444 avss.n584 avss.n542 8.61832
R1445 avss.n585 avss.n584 8.61832
R1446 avss.n586 avss.n540 8.61832
R1447 avss.n593 avss.n540 8.61832
R1448 avss.n535 avss.n527 8.61832
R1449 avss.n603 avss.n535 8.61832
R1450 avss.n603 avss.n602 8.61832
R1451 avss.n601 avss.n536 8.61832
R1452 avss.n595 avss.n536 8.61832
R1453 avss.n595 avss.n594 8.61832
R1454 avss.n561 avss.n560 8.61832
R1455 avss.n560 avss.n559 8.61832
R1456 avss.n554 avss.n526 8.61832
R1457 avss.t159 avss.t316 8.6067
R1458 avss.n672 avss.n671 8.4666
R1459 avss.n667 avss.n338 8.37766
R1460 avss.n347 avss.n338 8.37766
R1461 avss.n727 avss.n310 8.11041
R1462 avss.n727 avss.n726 8.11041
R1463 avss.n330 avss.n294 8.02619
R1464 avss.n671 avss.n330 8.00675
R1465 avss.t215 avss.t170 7.9692
R1466 avss.n347 avss.n337 7.938
R1467 avss.n667 avss.n337 7.938
R1468 avss.n334 avss.n333 7.48375
R1469 avss.n499 avss.n496 7.46717
R1470 avss.n501 avss.n500 7.46717
R1471 avss.n492 avss.n490 7.46717
R1472 avss.n487 avss.n478 7.46717
R1473 avss.n619 avss.n476 7.19646
R1474 avss.n670 avss.n334 7.16066
R1475 avss.t57 avss.t2 7.01296
R1476 avss.n333 avss.n329 6.89147
R1477 avss.n329 avss.n294 6.89083
R1478 avss.n308 avss.n306 6.88285
R1479 avss.n395 avss.n308 6.88285
R1480 avss.n309 avss.n307 6.88285
R1481 avss.n679 avss.n309 6.88285
R1482 avss.n341 avss.n339 6.5005
R1483 avss.t70 avss.n341 6.5005
R1484 avss.n342 avss.n340 6.5005
R1485 avss.t70 avss.n342 6.5005
R1486 avss.n442 avss.n387 6.48963
R1487 avss.n641 avss.n368 6.47706
R1488 avss.n641 avss.n639 6.47706
R1489 avss.n647 avss.n365 6.47706
R1490 avss.n647 avss.n366 6.47706
R1491 avss.n610 avss.n526 6.46387
R1492 avss.n618 avss.n293 6.2535
R1493 avss.n770 avss.n6 6.05765
R1494 avss.t175 avss.t176 6.05672
R1495 avss.n729 avss.n728 5.90959
R1496 avss.n730 avss.n729 5.90959
R1497 avss.n732 avss.n731 5.90959
R1498 avss.n731 avss.n730 5.90959
R1499 avss.n443 avss.n442 5.79451
R1500 avss.n771 avss.n770 5.78505
R1501 avss.n669 avss.n668 5.7846
R1502 avss.n336 avss.n335 5.76099
R1503 avss.n345 avss.n344 5.76099
R1504 avss.n305 avss.n304 5.70305
R1505 avss.n699 avss.n698 5.70305
R1506 avss.n712 avss.n711 5.70305
R1507 avss.n714 avss.n713 5.70305
R1508 avss.n312 avss.n310 5.70305
R1509 avss.n347 avss.n346 5.6605
R1510 avss.n297 avss.n296 5.6605
R1511 avss.n304 avss.n303 5.6605
R1512 avss.n735 avss.n734 5.6605
R1513 avss.n692 avss.n691 5.6605
R1514 avss.n698 avss.n697 5.6605
R1515 avss.n690 avss.n298 5.6605
R1516 avss.n705 avss.n704 5.6605
R1517 avss.n711 avss.n710 5.6605
R1518 avss.n703 avss.n702 5.6605
R1519 avss.n721 avss.n720 5.6605
R1520 avss.n715 avss.n714 5.6605
R1521 avss.n722 avss.n311 5.6605
R1522 avss.n319 avss.n318 5.6605
R1523 avss.n313 avss.n312 5.6605
R1524 avss.n726 avss.n725 5.6605
R1525 avss.n668 avss.n667 5.6605
R1526 avss.n433 avss.n391 5.27077
R1527 avss.n437 avss.n391 5.27077
R1528 avss.n428 avss.n390 5.27077
R1529 avss.n437 avss.n390 5.27077
R1530 avss.n331 avss.n326 5.27077
R1531 avss.n354 avss.n326 5.27077
R1532 avss.n674 avss.n327 5.27077
R1533 avss.n352 avss.n327 5.27077
R1534 avss.n636 avss.n366 5.07277
R1535 avss.n647 avss.n646 5.07277
R1536 avss.n460 avss.n365 5.07277
R1537 avss.n440 avss.n439 5.0436
R1538 avss.n439 avss.n438 5.0436
R1539 avss.n435 avss.n434 5.0436
R1540 avss.n673 avss.n332 5.0436
R1541 avss.n351 avss.n332 5.0436
R1542 avss.n677 avss.n676 5.0436
R1543 avss.n678 avss.n677 5.0436
R1544 avss.n522 avss.n521 5.0005
R1545 avss.n521 avss.n520 5.0005
R1546 avss.n513 avss.n509 5.0005
R1547 avss.n519 avss.n513 5.0005
R1548 avss.n517 avss.n516 5.0005
R1549 avss.n518 avss.n517 5.0005
R1550 avss.n515 avss.n512 5.0005
R1551 avss.n514 avss.n512 5.0005
R1552 avss.n639 avss.n638 4.95167
R1553 avss.n461 avss.n368 4.95167
R1554 avss.n740 avss.n17 4.86769
R1555 avss.n24 avss.n22 4.6805
R1556 avss.t85 avss.n24 4.6805
R1557 avss.n272 avss.n25 4.6805
R1558 avss.t85 avss.n25 4.6805
R1559 avss.n630 avss.n629 4.5005
R1560 avss.n632 avss.n631 4.5005
R1561 avss.n642 avss.n641 4.5005
R1562 avss.n634 avss.n633 4.5005
R1563 avss.n628 avss.n369 4.5005
R1564 avss.n458 avss.n371 4.5005
R1565 avss.n464 avss.n463 4.5005
R1566 avss.n468 avss.n467 4.5005
R1567 avss.n466 avss.n465 4.5005
R1568 avss.n510 avss.n507 4.3603
R1569 avss.n524 avss.n508 4.34678
R1570 avss.n510 avss.n508 4.34003
R1571 avss.n442 avss.n386 4.22604
R1572 avss.n620 avss.n619 4.21323
R1573 avss.n754 avss.n18 4.04961
R1574 avss.n346 avss.n320 4.00655
R1575 avss.n648 avss.n361 3.9532
R1576 avss.n448 avss.n361 3.9532
R1577 avss.n640 avss.n360 3.9532
R1578 avss.n448 avss.n360 3.9532
R1579 avss.n770 avss.n769 3.94537
R1580 avss.t366 avss.t264 3.7849
R1581 avss.n525 avss.n524 3.78259
R1582 avss.n465 avss.n457 3.77378
R1583 avss.n642 avss.n367 3.77209
R1584 avss.n633 avss.n370 3.77014
R1585 avss.n688 avss.n687 3.68964
R1586 avss.n736 avss.n735 3.57087
R1587 avss.n690 avss.n295 3.57087
R1588 avss.n703 avss.n689 3.57087
R1589 avss.n723 avss.n722 3.57087
R1590 avss.n725 avss.n724 3.57087
R1591 avss.n616 avss.n615 3.4105
R1592 avss.n381 avss.n380 3.4105
R1593 avss.n299 avss.t289 3.3065
R1594 avss.n299 avss.t111 3.3065
R1595 avss.t89 avss.n302 3.3065
R1596 avss.n302 avss.t288 3.3065
R1597 avss.n693 avss.t293 3.3065
R1598 avss.n693 avss.t102 3.3065
R1599 avss.t118 avss.n696 3.3065
R1600 avss.n696 avss.t290 3.3065
R1601 avss.n706 avss.t286 3.3065
R1602 avss.n706 avss.t143 3.3065
R1603 avss.t62 avss.n709 3.3065
R1604 avss.n709 avss.t284 3.3065
R1605 avss.n718 avss.t291 3.3065
R1606 avss.n718 avss.t140 3.3065
R1607 avss.n716 avss.t146 3.3065
R1608 avss.n716 avss.t294 3.3065
R1609 avss.n316 avss.t287 3.3065
R1610 avss.n316 avss.t73 3.3065
R1611 avss.n314 avss.t94 3.3065
R1612 avss.n314 avss.t292 3.3065
R1613 avss.n412 avss.t3 3.3065
R1614 avss.n412 avss.t1 3.3065
R1615 avss.n466 avss.n368 3.23878
R1616 avss.n639 avss.n634 3.23878
R1617 avss.n467 avss.n365 3.23878
R1618 avss.n369 avss.n366 3.23878
R1619 avss.t72 avss.t175 3.18798
R1620 avss.n611 avss.n610 3.1005
R1621 avss.n768 avss.n7 2.6005
R1622 avss.t200 avss.t340 2.52344
R1623 avss.n726 avss.n311 2.42291
R1624 avss.n702 avss.n311 2.42291
R1625 avss.n734 avss.n298 2.42291
R1626 avss.n699 avss.n305 2.42291
R1627 avss.n713 avss.n712 2.42291
R1628 avss.n713 avss.n310 2.42291
R1629 avss.n577 avss.n542 2.40842
R1630 avss.n594 avss.n593 2.40842
R1631 avss.n612 avss.n506 2.32925
R1632 avss.n737 avss.n294 2.31886
R1633 avss.n333 avss.n320 2.31886
R1634 avss.n561 avss.n550 2.28169
R1635 avss.n609 avss.n527 2.28169
R1636 avss.n515 avss.n511 2.25932
R1637 avss.n670 avss.n669 2.2505
R1638 avss.n754 avss.n753 2.2505
R1639 avss.n611 avss.n525 2.17339
R1640 avss.n610 avss.n609 2.15496
R1641 avss.n619 avss.n618 2.1358
R1642 avss.n467 avss.n466 2.11769
R1643 avss.n634 avss.n369 2.11769
R1644 avss.n738 avss.n293 2.058
R1645 avss.n267 avss.t4 1.99563
R1646 avss.t298 avss.n268 1.8927
R1647 avss.n617 avss.n616 1.80585
R1648 avss.n701 avss.n298 1.80222
R1649 avss.n700 avss.n699 1.80222
R1650 avss.n275 avss.n274 1.6605
R1651 avss.n730 avss.t320 1.59424
R1652 avss.n370 avss.n367 1.58008
R1653 avss.n457 avss.n367 1.58008
R1654 avss.n751 avss.n20 1.48467
R1655 avss.n618 avss.n617 1.40612
R1656 avss.n292 avss.n291 1.34141
R1657 avss.n274 avss.n19 1.338
R1658 avss.n750 avss.n21 1.32209
R1659 avss.n741 avss.n276 1.27675
R1660 avss.n279 avss.n278 1.14936
R1661 avss.n287 avss.n286 1.14936
R1662 avss.n286 avss.n285 1.14839
R1663 avss.n278 avss.n277 1.14811
R1664 avss.n277 avss.n21 1.08686
R1665 avss.n280 avss.n279 1.08686
R1666 avss.n281 avss.n280 1.08686
R1667 avss.n283 avss.n282 1.08686
R1668 avss.n288 avss.n287 1.08686
R1669 avss.n289 avss.n288 1.08686
R1670 avss.n290 avss.n289 1.08686
R1671 avss.n291 avss.n290 1.08686
R1672 avss.n282 avss.n281 1.08005
R1673 avss.n301 avss.n300 1.05355
R1674 avss.n695 avss.n694 1.05355
R1675 avss.n708 avss.n707 1.05355
R1676 avss.n719 avss.n717 1.05355
R1677 avss.n317 avss.n315 1.05355
R1678 avss.n276 avss.n275 1.00987
R1679 avss.n285 avss.n284 1.00505
R1680 avss.n761 avss.n760 1.00393
R1681 avss.t48 avss.n761 1.00393
R1682 avss.n755 avss.n12 1.00393
R1683 avss.t48 avss.n12 1.00393
R1684 avss.t225 avss.t167 0.956745
R1685 avss.n343 avss.n336 0.955426
R1686 avss.n345 avss.n343 0.953203
R1687 avss.n739 avss.n292 0.902375
R1688 avss.n752 avss.n751 0.839875
R1689 avss.n153 avss.n6 0.79175
R1690 avss.n523 avss.n509 0.753441
R1691 avss.n379 avss.n377 0.695812
R1692 avss.n632 avss.n630 0.695812
R1693 avss.n638 avss.n636 0.695812
R1694 avss.n646 avss.n644 0.695812
R1695 avss.n461 avss.n460 0.695812
R1696 avss.n464 avss.n371 0.695812
R1697 avss.n614 avss.n613 0.695812
R1698 avss.n375 avss.n373 0.679185
R1699 avss.n380 avss.n379 0.654797
R1700 avss.t61 avss.n419 0.637996
R1701 avss.n687 avss.n321 0.635318
R1702 avss.n702 avss.n701 0.62119
R1703 avss.n712 avss.n700 0.62119
R1704 avss.n630 avss.n628 0.572766
R1705 avss.n468 avss.n371 0.572766
R1706 avss.n525 avss.n507 0.571446
R1707 avss.n304 avss.n301 0.527027
R1708 avss.n300 avss.n297 0.527027
R1709 avss.n698 avss.n695 0.527027
R1710 avss.n694 avss.n692 0.527027
R1711 avss.n711 avss.n708 0.527027
R1712 avss.n707 avss.n705 0.527027
R1713 avss.n717 avss.n714 0.527027
R1714 avss.n721 avss.n719 0.527027
R1715 avss.n315 avss.n312 0.527027
R1716 avss.n319 avss.n317 0.527027
R1717 avss.n688 avss.n320 0.505881
R1718 avss.n724 avss.n688 0.497189
R1719 avss.n724 avss.n723 0.478977
R1720 avss.n723 avss.n689 0.478977
R1721 avss.n689 avss.n295 0.478977
R1722 avss.n736 avss.n295 0.478977
R1723 avss.n627 avss.n626 0.46925
R1724 avss.n626 avss.n625 0.46925
R1725 avss.n625 avss.n624 0.46925
R1726 avss.n624 avss.n623 0.46925
R1727 avss.n623 avss.n622 0.46925
R1728 avss.n622 avss.n621 0.46925
R1729 avss.n621 avss.n620 0.46925
R1730 avss.n470 avss.n469 0.46925
R1731 avss.n471 avss.n470 0.46925
R1732 avss.n472 avss.n471 0.46925
R1733 avss.n473 avss.n472 0.46925
R1734 avss.n474 avss.n473 0.46925
R1735 avss.n475 avss.n474 0.46925
R1736 avss.n476 avss.n475 0.46925
R1737 avss.n633 avss.n632 0.451672
R1738 avss.n644 avss.n642 0.451672
R1739 avss.n465 avss.n464 0.451672
R1740 avss.n738 avss.n737 0.387296
R1741 avss.n737 avss.n736 0.380881
R1742 avss.n292 avss.n6 0.364875
R1743 avss.n351 avss.t341 0.319248
R1744 avss.n615 avss.n614 0.311047
R1745 avss.n414 avss.n413 0.291392
R1746 avss.n413 avss.n411 0.291392
R1747 avss.n511 avss.n510 0.274029
R1748 avss.n522 avss.n508 0.266214
R1749 avss.n524 avss.n523 0.266214
R1750 avss.n516 avss.n507 0.266214
R1751 avss.n256 avss 0.248811
R1752 avss avss.n251 0.248811
R1753 avss.n242 avss 0.248811
R1754 avss avss.n237 0.248811
R1755 avss.n228 avss 0.248811
R1756 avss avss.n223 0.248811
R1757 avss.n214 avss 0.248811
R1758 avss avss.n209 0.248811
R1759 avss.n200 avss 0.248811
R1760 avss avss.n195 0.248811
R1761 avss.n186 avss 0.248811
R1762 avss avss.n181 0.248811
R1763 avss.n172 avss 0.248811
R1764 avss avss.n167 0.248811
R1765 avss.n158 avss 0.248811
R1766 avss.n616 avss.n370 0.237405
R1767 avss.n388 avss.n386 0.216779
R1768 avss.n403 avss.n402 0.182466
R1769 avss.n752 avss.n19 0.153
R1770 avss.n757 avss.n16 0.152959
R1771 avss.n18 avss.n15 0.152959
R1772 avss.n389 avss.n387 0.141409
R1773 avss.n751 avss.n750 0.128909
R1774 avss.n415 avss.n400 0.119588
R1775 avss.n457 avss.n456 0.118318
R1776 avss.n701 avss.n307 0.11675
R1777 avss.n700 avss.n306 0.11675
R1778 avss.n402 avss.n401 0.11673
R1779 avss.n456 avss.n381 0.114189
R1780 avss.n401 avss.n321 0.113554
R1781 avss.n339 avss.n337 0.109912
R1782 avss.n340 avss.n338 0.109912
R1783 avss avss.n153 0.107764
R1784 avss.n740 avss.n739 0.10175
R1785 avss.n728 avss.n727 0.0994362
R1786 avss.n733 avss.n732 0.0994362
R1787 avss.n430 avss.n429 0.0907913
R1788 avss.n334 avss.n331 0.0890714
R1789 avss.n674 avss.n330 0.0890714
R1790 avss.n433 avss.n432 0.0890714
R1791 avss.n676 avss.n329 0.0866111
R1792 avss.n673 avss.n672 0.0850455
R1793 avss.n434 avss.n431 0.0850455
R1794 avss.n284 avss.n283 0.0823182
R1795 avss.n28 avss.n20 0.0815811
R1796 avss.n256 avss.n255 0.0815811
R1797 avss.n251 avss.n37 0.0815811
R1798 avss.n242 avss.n241 0.0815811
R1799 avss.n237 avss.n53 0.0815811
R1800 avss.n228 avss.n227 0.0815811
R1801 avss.n223 avss.n69 0.0815811
R1802 avss.n214 avss.n213 0.0815811
R1803 avss.n209 avss.n85 0.0815811
R1804 avss.n200 avss.n199 0.0815811
R1805 avss.n195 avss.n101 0.0815811
R1806 avss.n186 avss.n185 0.0815811
R1807 avss.n181 avss.n117 0.0815811
R1808 avss.n172 avss.n171 0.0815811
R1809 avss.n167 avss.n133 0.0815811
R1810 avss.n158 avss.n157 0.0815811
R1811 avss.n778 avss.n0 0.0815811
R1812 avss.n284 avss.n269 0.0793136
R1813 avss.n612 avss.n611 0.0784703
R1814 avss.n641 avss.n640 0.0674065
R1815 avss.n648 avss.n647 0.0674065
R1816 avss.n33 avss.n29 0.0553986
R1817 avss.n254 avss.n36 0.0553986
R1818 avss.n49 avss.n48 0.0553986
R1819 avss.n240 avss.n52 0.0553986
R1820 avss.n65 avss.n64 0.0553986
R1821 avss.n226 avss.n68 0.0553986
R1822 avss.n81 avss.n80 0.0553986
R1823 avss.n212 avss.n84 0.0553986
R1824 avss.n97 avss.n96 0.0553986
R1825 avss.n198 avss.n100 0.0553986
R1826 avss.n113 avss.n112 0.0553986
R1827 avss.n184 avss.n116 0.0553986
R1828 avss.n129 avss.n128 0.0553986
R1829 avss.n170 avss.n132 0.0553986
R1830 avss.n145 avss.n144 0.0553986
R1831 avss.n156 avss.n152 0.0553986
R1832 avss.n410 avss.n403 0.0538514
R1833 avss.n443 avss.n381 0.0532162
R1834 avss.n153 avss 0.04675
R1835 avss.n668 avss.n336 0.0436892
R1836 avss.n735 avss.n297 0.0430541
R1837 avss.n692 avss.n690 0.0430541
R1838 avss.n705 avss.n703 0.0430541
R1839 avss.n722 avss.n721 0.0430541
R1840 avss.n725 avss.n319 0.0430541
R1841 avss.n415 avss.n414 0.0430541
R1842 avss.n346 avss.n345 0.0430541
R1843 avss.n411 avss.n410 0.0427365
R1844 avss avss.n778 0.0410405
R1845 avss avss.n35 0.0351284
R1846 avss.n252 avss 0.0351284
R1847 avss avss.n51 0.0351284
R1848 avss.n238 avss 0.0351284
R1849 avss avss.n67 0.0351284
R1850 avss.n224 avss 0.0351284
R1851 avss avss.n83 0.0351284
R1852 avss.n210 avss 0.0351284
R1853 avss avss.n99 0.0351284
R1854 avss.n196 avss 0.0351284
R1855 avss avss.n115 0.0351284
R1856 avss.n182 avss 0.0351284
R1857 avss avss.n131 0.0351284
R1858 avss.n168 avss 0.0351284
R1859 avss avss.n147 0.0351284
R1860 avss.n154 avss 0.0351284
R1861 avss.n771 avss.n5 0.0334392
R1862 avss.n33 avss.n28 0.0266824
R1863 avss.n255 avss.n254 0.0266824
R1864 avss.n49 avss.n37 0.0266824
R1865 avss.n241 avss.n240 0.0266824
R1866 avss.n65 avss.n53 0.0266824
R1867 avss.n227 avss.n226 0.0266824
R1868 avss.n81 avss.n69 0.0266824
R1869 avss.n213 avss.n212 0.0266824
R1870 avss.n97 avss.n85 0.0266824
R1871 avss.n199 avss.n198 0.0266824
R1872 avss.n113 avss.n101 0.0266824
R1873 avss.n185 avss.n184 0.0266824
R1874 avss.n129 avss.n117 0.0266824
R1875 avss.n171 avss.n170 0.0266824
R1876 avss.n145 avss.n133 0.0266824
R1877 avss.n157 avss.n156 0.0266824
R1878 avss.n5 avss.n0 0.0266824
R1879 avss.n772 avss.n771 0.0224595
R1880 avss.n380 avss.n375 0.0190811
R1881 avss.n756 avss.n755 0.0173784
R1882 avss.n759 avss.n758 0.0173478
R1883 avss.n35 avss.n29 0.00641216
R1884 avss.n252 avss.n36 0.00641216
R1885 avss.n51 avss.n48 0.00641216
R1886 avss.n238 avss.n52 0.00641216
R1887 avss.n67 avss.n64 0.00641216
R1888 avss.n224 avss.n68 0.00641216
R1889 avss.n83 avss.n80 0.00641216
R1890 avss.n210 avss.n84 0.00641216
R1891 avss.n99 avss.n96 0.00641216
R1892 avss.n196 avss.n100 0.00641216
R1893 avss.n115 avss.n112 0.00641216
R1894 avss.n182 avss.n116 0.00641216
R1895 avss.n131 avss.n128 0.00641216
R1896 avss.n168 avss.n132 0.00641216
R1897 avss.n147 avss.n144 0.00641216
R1898 avss.n154 avss.n152 0.00641216
R1899 avss.n741 avss.n740 0.004875
R1900 dvss.n905 dvss.n903 198880
R1901 dvss.n905 dvss.t259 192115
R1902 dvss.n2668 dvss.n2667 39445.1
R1903 dvss.n902 dvss.n900 33375.3
R1904 dvss.n58 dvss.n14 22266.3
R1905 dvss.n856 dvss.n855 9262.6
R1906 dvss.n3641 dvss.n120 8941.81
R1907 dvss.n676 dvss.t131 8003.11
R1908 dvss.t483 dvss.n146 8003.11
R1909 dvss.t448 dvss.n296 8003.11
R1910 dvss.t530 dvss.n2671 8003.11
R1911 dvss.t360 dvss.n360 8003.11
R1912 dvss.t283 dvss.n1806 8003.11
R1913 dvss.n1513 dvss.t195 8003.11
R1914 dvss.t222 dvss.n1226 8003.11
R1915 dvss.n1004 dvss.t38 8003.11
R1916 dvss.n14 dvss.n13 7873.38
R1917 dvss.t127 dvss.t125 7626.67
R1918 dvss.t133 dvss.t131 7626.67
R1919 dvss.t479 dvss.t477 7626.67
R1920 dvss.t483 dvss.t481 7626.67
R1921 dvss.t444 dvss.t442 7626.67
R1922 dvss.t448 dvss.t446 7626.67
R1923 dvss.t526 dvss.t524 7626.67
R1924 dvss.t530 dvss.t528 7626.67
R1925 dvss.t356 dvss.t354 7626.67
R1926 dvss.t360 dvss.t358 7626.67
R1927 dvss.t287 dvss.t291 7626.67
R1928 dvss.t283 dvss.t285 7626.67
R1929 dvss.t197 dvss.t199 7626.67
R1930 dvss.t203 dvss.t195 7626.67
R1931 dvss.t216 dvss.t218 7626.67
R1932 dvss.t222 dvss.t214 7626.67
R1933 dvss.t36 dvss.t40 7626.67
R1934 dvss.t44 dvss.t38 7626.67
R1935 dvss.n3571 dvss.n162 6332.05
R1936 dvss.n1849 dvss.n1784 6332.05
R1937 dvss.n1879 dvss.n1878 6332.05
R1938 dvss.n1824 dvss.n1790 6332.05
R1939 dvss.n1796 dvss.n1795 6332.05
R1940 dvss.n1594 dvss.n494 6332.05
R1941 dvss.n1216 dvss.n1215 6332.05
R1942 dvss.n1121 dvss.n604 6332.05
R1943 dvss.n1292 dvss.t78 6153.5
R1944 dvss.n2882 dvss.t78 6153.5
R1945 dvss.t97 dvss.n134 6153.5
R1946 dvss.n3547 dvss.t493 6153.5
R1947 dvss.t78 dvss.n398 6153.5
R1948 dvss.n1581 dvss.t78 6153.5
R1949 dvss.n1108 dvss.t78 6153.5
R1950 dvss.n3651 dvss.n3650 5772.37
R1951 dvss.n3650 dvss.n120 5605.26
R1952 dvss.n58 dvss 5162.25
R1953 dvss.n3636 dvss.n134 5082
R1954 dvss.n1871 dvss.n272 5082
R1955 dvss.n3548 dvss.n3547 5082
R1956 dvss.n2224 dvss.n336 5082
R1957 dvss.n2272 dvss.n272 5082
R1958 dvss.n1846 dvss.n336 5082
R1959 dvss.n1821 dvss.n398 5082
R1960 dvss.n2882 dvss.n2881 5082
R1961 dvss.n1582 dvss.n1581 5082
R1962 dvss.n1292 dvss.n1291 5082
R1963 dvss.n1109 dvss.n1108 5082
R1964 dvss.t261 dvss.n903 4455
R1965 dvss.n61 dvss.n11 4160.18
R1966 dvss.n61 dvss.n12 4160.18
R1967 dvss.n62 dvss.n11 4160.18
R1968 dvss.n62 dvss.n12 4160.18
R1969 dvss.t177 dvss.n14 3236.46
R1970 dvss.t259 dvss.t261 2310
R1971 dvss.t99 dvss.t93 1778.24
R1972 dvss.t487 dvss.t495 1778.24
R1973 dvss.t99 dvss.n146 1652.85
R1974 dvss.n2671 dvss.t487 1652.85
R1975 dvss.n13 dvss.t380 1124.77
R1976 dvss.t111 dvss.n59 1124.77
R1977 dvss.n2667 dvss.t78 1094.3
R1978 dvss.n863 dvss.n856 1069.72
R1979 dvss.n860 dvss.n859 1013.99
R1980 dvss.n59 dvss.n58 996.557
R1981 dvss.t380 dvss.t429 920.795
R1982 dvss.t344 dvss.t429 920.795
R1983 dvss.t344 dvss.t113 920.795
R1984 dvss.t113 dvss.t111 920.795
R1985 dvss.n855 dvss.n854 769.572
R1986 dvss.n3642 dvss.n3641 769.572
R1987 dvss.n861 dvss.n860 769.572
R1988 dvss.t60 dvss.n146 761.905
R1989 dvss.n2671 dvss.t34 761.905
R1990 dvss.t22 dvss.n296 761.905
R1991 dvss.t12 dvss.n360 761.905
R1992 dvss.n1806 dvss.t272 761.905
R1993 dvss.n1513 dvss.t366 761.905
R1994 dvss.n1226 dvss.t461 761.905
R1995 dvss.n676 dvss.t238 761.905
R1996 dvss.n1004 dvss.t68 761.905
R1997 dvss.n3438 dvss.n3437 747.437
R1998 dvss.n3254 dvss.n269 747.437
R1999 dvss.n3138 dvss.n333 747.437
R2000 dvss.n3035 dvss.n391 747.437
R2001 dvss.n2915 dvss.n448 747.437
R2002 dvss.n1488 dvss.n1476 747.437
R2003 dvss.n1323 dvss.n557 747.437
R2004 dvss.n1100 dvss.n1099 747.437
R2005 dvss.n1889 dvss.n85 607.51
R2006 dvss.n176 dvss.n113 607.51
R2007 dvss.n1890 dvss.n84 592.001
R2008 dvss.n177 dvss.n112 592.001
R2009 dvss.n3573 dvss.n156 590.068
R2010 dvss.n1853 dvss.n1852 590.068
R2011 dvss.n1883 dvss.n1882 590.068
R2012 dvss.n1828 dvss.n1827 590.068
R2013 dvss.n1801 dvss.n1800 590.068
R2014 dvss.n1608 dvss.n1607 590.068
R2015 dvss.n1221 dvss.n1220 590.068
R2016 dvss.n1135 dvss.n1134 590.068
R2017 dvss.n848 dvss.n772 590.068
R2018 dvss.n1891 dvss.n1888 588.516
R2019 dvss.n178 dvss.n171 588.516
R2020 dvss.n3592 dvss.n3591 587.271
R2021 dvss.n1856 dvss.n1779 587.271
R2022 dvss.n1886 dvss.n1778 587.271
R2023 dvss.n1831 dvss.n1785 587.271
R2024 dvss.n1804 dvss.n1791 587.271
R2025 dvss.n1621 dvss.n485 587.271
R2026 dvss.n1224 dvss.n1211 587.271
R2027 dvss.n1148 dvss.n595 587.271
R2028 dvss.n842 dvss.n841 587.271
R2029 dvss.n1319 dvss.n561 585
R2030 dvss.n561 dvss.n557 585
R2031 dvss.n1310 dvss.n564 585
R2032 dvss.n1313 dvss.n1312 585
R2033 dvss.n1309 dvss.n553 585
R2034 dvss.n1309 dvss.n557 585
R2035 dvss.n551 dvss.n550 585
R2036 dvss.n1324 dvss.n550 585
R2037 dvss.n1336 dvss.n1335 585
R2038 dvss.n1337 dvss.n1336 585
R2039 dvss.n547 dvss.n546 585
R2040 dvss.n1338 dvss.n546 585
R2041 dvss.n1349 dvss.n1348 585
R2042 dvss.n1349 dvss.n544 585
R2043 dvss.n1350 dvss.n539 585
R2044 dvss.n1351 dvss.n1350 585
R2045 dvss.n1363 dvss.n540 585
R2046 dvss.n545 dvss.n540 585
R2047 dvss.n1364 dvss.n535 585
R2048 dvss.n1369 dvss.n535 585
R2049 dvss.n1373 dvss.n536 585
R2050 dvss.n1373 dvss.n1372 585
R2051 dvss.n1374 dvss.n530 585
R2052 dvss.n1375 dvss.n1374 585
R2053 dvss.n1384 dvss.n531 585
R2054 dvss.n1225 dvss.n531 585
R2055 dvss.n1385 dvss.n525 585
R2056 dvss.n527 dvss.n525 585
R2057 dvss.n1398 dvss.n526 585
R2058 dvss.n1398 dvss.n1397 585
R2059 dvss.n1399 dvss.n518 585
R2060 dvss.n1400 dvss.n1399 585
R2061 dvss.n524 dvss.n523 585
R2062 dvss.n1401 dvss.n524 585
R2063 dvss.n1405 dvss.n1404 585
R2064 dvss.n1404 dvss.n1403 585
R2065 dvss.n509 dvss.n507 585
R2066 dvss.n507 dvss.n504 585
R2067 dvss.n1579 dvss.n1578 585
R2068 dvss.n1580 dvss.n1579 585
R2069 dvss.n510 dvss.n508 585
R2070 dvss.n508 dvss.n506 585
R2071 dvss.n1486 dvss.n1420 585
R2072 dvss.n1485 dvss.n1421 585
R2073 dvss.n1484 dvss.n1425 585
R2074 dvss.n1490 dvss.n1426 585
R2075 dvss.n1492 dvss.n1491 585
R2076 dvss.n1493 dvss.n1492 585
R2077 dvss.n1475 dvss.n1430 585
R2078 dvss.n1494 dvss.n1475 585
R2079 dvss.n1496 dvss.n1435 585
R2080 dvss.n1496 dvss.n1495 585
R2081 dvss.n1498 dvss.n1497 585
R2082 dvss.n1497 dvss.n1472 585
R2083 dvss.n1502 dvss.n1501 585
R2084 dvss.n1503 dvss.n1502 585
R2085 dvss.n1471 dvss.n1441 585
R2086 dvss.n1504 dvss.n1471 585
R2087 dvss.n1507 dvss.n1446 585
R2088 dvss.n1507 dvss.n1506 585
R2089 dvss.n1508 dvss.n1447 585
R2090 dvss.n1509 dvss.n1508 585
R2091 dvss.n1469 dvss.n1468 585
R2092 dvss.n1512 dvss.n1469 585
R2093 dvss.n1515 dvss.n1450 585
R2094 dvss.n1515 dvss.n1514 585
R2095 dvss.n1516 dvss.n1458 585
R2096 dvss.n1517 dvss.n1516 585
R2097 dvss.n1466 dvss.n1459 585
R2098 dvss.n1518 dvss.n1466 585
R2099 dvss.n1522 dvss.n1467 585
R2100 dvss.n1522 dvss.n1521 585
R2101 dvss.n1523 dvss.n1463 585
R2102 dvss.n1524 dvss.n1523 585
R2103 dvss.n459 dvss.n458 585
R2104 dvss.n1525 dvss.n459 585
R2105 dvss.n2885 dvss.n2884 585
R2106 dvss.n2884 dvss.n2883 585
R2107 dvss.n453 dvss.n451 585
R2108 dvss.n451 dvss.n449 585
R2109 dvss.n2913 dvss.n2912 585
R2110 dvss.n2914 dvss.n2913 585
R2111 dvss.n454 dvss.n452 585
R2112 dvss.n2901 dvss.n2899 585
R2113 dvss.n2905 dvss.n2904 585
R2114 dvss.n2902 dvss.n444 585
R2115 dvss.n442 dvss.n441 585
R2116 dvss.n2916 dvss.n441 585
R2117 dvss.n2928 dvss.n2927 585
R2118 dvss.n2929 dvss.n2928 585
R2119 dvss.n438 dvss.n437 585
R2120 dvss.n2930 dvss.n437 585
R2121 dvss.n2941 dvss.n2940 585
R2122 dvss.n2941 dvss.n435 585
R2123 dvss.n2942 dvss.n430 585
R2124 dvss.n2943 dvss.n2942 585
R2125 dvss.n2955 dvss.n431 585
R2126 dvss.n436 dvss.n431 585
R2127 dvss.n2956 dvss.n426 585
R2128 dvss.n2961 dvss.n426 585
R2129 dvss.n2965 dvss.n427 585
R2130 dvss.n2965 dvss.n2964 585
R2131 dvss.n2966 dvss.n421 585
R2132 dvss.n2967 dvss.n2966 585
R2133 dvss.n2976 dvss.n422 585
R2134 dvss.n1805 dvss.n422 585
R2135 dvss.n2977 dvss.n416 585
R2136 dvss.n418 dvss.n416 585
R2137 dvss.n2990 dvss.n417 585
R2138 dvss.n2990 dvss.n2989 585
R2139 dvss.n2991 dvss.n409 585
R2140 dvss.n2992 dvss.n2991 585
R2141 dvss.n415 dvss.n414 585
R2142 dvss.n2993 dvss.n415 585
R2143 dvss.n2998 dvss.n2997 585
R2144 dvss.n2997 dvss.n2996 585
R2145 dvss.n400 dvss.n399 585
R2146 dvss.n2995 dvss.n399 585
R2147 dvss.n3014 dvss.n3013 585
R2148 dvss.n3015 dvss.n3014 585
R2149 dvss.n394 dvss.n393 585
R2150 dvss.n3016 dvss.n393 585
R2151 dvss.n3033 dvss.n3032 585
R2152 dvss.n395 dvss.n392 585
R2153 dvss.n389 dvss.n388 585
R2154 dvss.n3038 dvss.n3037 585
R2155 dvss.n383 dvss.n382 585
R2156 dvss.n390 dvss.n382 585
R2157 dvss.n3050 dvss.n3049 585
R2158 dvss.n3051 dvss.n3050 585
R2159 dvss.n379 dvss.n378 585
R2160 dvss.n3052 dvss.n379 585
R2161 dvss.n3058 dvss.n3057 585
R2162 dvss.n3057 dvss.n3056 585
R2163 dvss.n373 dvss.n372 585
R2164 dvss.n3055 dvss.n372 585
R2165 dvss.n3076 dvss.n3075 585
R2166 dvss.n3077 dvss.n3076 585
R2167 dvss.n367 dvss.n366 585
R2168 dvss.n369 dvss.n367 585
R2169 dvss.n3082 dvss.n3081 585
R2170 dvss.n3081 dvss.n3080 585
R2171 dvss.n362 dvss.n361 585
R2172 dvss.n368 dvss.n361 585
R2173 dvss.n3093 dvss.n3092 585
R2174 dvss.n3094 dvss.n3093 585
R2175 dvss.n357 dvss.n356 585
R2176 dvss.n356 dvss.n354 585
R2177 dvss.n3107 dvss.n3106 585
R2178 dvss.n3108 dvss.n3107 585
R2179 dvss.n352 dvss.n346 585
R2180 dvss.n3109 dvss.n352 585
R2181 dvss.n3115 dvss.n3114 585
R2182 dvss.n3114 dvss.n3113 585
R2183 dvss.n353 dvss.n340 585
R2184 dvss.n3112 dvss.n353 585
R2185 dvss.n3127 dvss.n341 585
R2186 dvss.n3111 dvss.n341 585
R2187 dvss.n3128 dvss.n334 585
R2188 dvss.n3133 dvss.n334 585
R2189 dvss.n3135 dvss.n335 585
R2190 dvss.n3135 dvss.n3134 585
R2191 dvss.n3136 dvss.n328 585
R2192 dvss.n330 dvss.n329 585
R2193 dvss.n3141 dvss.n3140 585
R2194 dvss.n331 dvss.n320 585
R2195 dvss.n318 dvss.n317 585
R2196 dvss.n332 dvss.n317 585
R2197 dvss.n3167 dvss.n3166 585
R2198 dvss.n3168 dvss.n3167 585
R2199 dvss.n314 dvss.n313 585
R2200 dvss.n3171 dvss.n314 585
R2201 dvss.n3175 dvss.n3174 585
R2202 dvss.n3174 dvss.n3173 585
R2203 dvss.n308 dvss.n307 585
R2204 dvss.n3172 dvss.n307 585
R2205 dvss.n3189 dvss.n3188 585
R2206 dvss.n3190 dvss.n3189 585
R2207 dvss.n303 dvss.n302 585
R2208 dvss.n3193 dvss.n303 585
R2209 dvss.n3198 dvss.n3197 585
R2210 dvss.n3197 dvss.n3196 585
R2211 dvss.n298 dvss.n297 585
R2212 dvss.n304 dvss.n297 585
R2213 dvss.n3209 dvss.n3208 585
R2214 dvss.n3210 dvss.n3209 585
R2215 dvss.n293 dvss.n292 585
R2216 dvss.n292 dvss.n290 585
R2217 dvss.n3223 dvss.n3222 585
R2218 dvss.n3224 dvss.n3223 585
R2219 dvss.n288 dvss.n282 585
R2220 dvss.n3225 dvss.n288 585
R2221 dvss.n3231 dvss.n3230 585
R2222 dvss.n3230 dvss.n3229 585
R2223 dvss.n289 dvss.n276 585
R2224 dvss.n3228 dvss.n289 585
R2225 dvss.n3243 dvss.n277 585
R2226 dvss.n3227 dvss.n277 585
R2227 dvss.n3244 dvss.n270 585
R2228 dvss.n3249 dvss.n270 585
R2229 dvss.n3251 dvss.n271 585
R2230 dvss.n3251 dvss.n3250 585
R2231 dvss.n3252 dvss.n264 585
R2232 dvss.n266 dvss.n265 585
R2233 dvss.n3257 dvss.n3256 585
R2234 dvss.n267 dvss.n255 585
R2235 dvss.n3275 dvss.n256 585
R2236 dvss.n268 dvss.n256 585
R2237 dvss.n3276 dvss.n251 585
R2238 dvss.n3286 dvss.n251 585
R2239 dvss.n3288 dvss.n252 585
R2240 dvss.n3288 dvss.n3287 585
R2241 dvss.n3289 dvss.n246 585
R2242 dvss.n3290 dvss.n3289 585
R2243 dvss.n241 dvss.n240 585
R2244 dvss.n250 dvss.n240 585
R2245 dvss.n3308 dvss.n3307 585
R2246 dvss.n3309 dvss.n3308 585
R2247 dvss.n242 dvss.n236 585
R2248 dvss.n238 dvss.n236 585
R2249 dvss.n3313 dvss.n237 585
R2250 dvss.n3313 dvss.n3312 585
R2251 dvss.n3314 dvss.n231 585
R2252 dvss.n3315 dvss.n3314 585
R2253 dvss.n3324 dvss.n232 585
R2254 dvss.n1887 dvss.n232 585
R2255 dvss.n3325 dvss.n226 585
R2256 dvss.n228 dvss.n226 585
R2257 dvss.n3338 dvss.n227 585
R2258 dvss.n3338 dvss.n3337 585
R2259 dvss.n3339 dvss.n219 585
R2260 dvss.n3340 dvss.n3339 585
R2261 dvss.n225 dvss.n224 585
R2262 dvss.n3341 dvss.n225 585
R2263 dvss.n3345 dvss.n3344 585
R2264 dvss.n3344 dvss.n3343 585
R2265 dvss.n210 dvss.n208 585
R2266 dvss.n208 dvss.n205 585
R2267 dvss.n3545 dvss.n3544 585
R2268 dvss.n3546 dvss.n3545 585
R2269 dvss.n211 dvss.n209 585
R2270 dvss.n209 dvss.n207 585
R2271 dvss.n3435 dvss.n3360 585
R2272 dvss.n3434 dvss.n3361 585
R2273 dvss.n3433 dvss.n3365 585
R2274 dvss.n3431 dvss.n3366 585
R2275 dvss.n3430 dvss.n3429 585
R2276 dvss.n3446 dvss.n3430 585
R2277 dvss.n3448 dvss.n3370 585
R2278 dvss.n3448 dvss.n3447 585
R2279 dvss.n3449 dvss.n3375 585
R2280 dvss.n3450 dvss.n3449 585
R2281 dvss.n3425 dvss.n3424 585
R2282 dvss.n3451 dvss.n3424 585
R2283 dvss.n3455 dvss.n3428 585
R2284 dvss.n3455 dvss.n3454 585
R2285 dvss.n3457 dvss.n3381 585
R2286 dvss.n3458 dvss.n3457 585
R2287 dvss.n3456 dvss.n3386 585
R2288 dvss.n3456 dvss.n3423 585
R2289 dvss.n3421 dvss.n3387 585
R2290 dvss.n3461 dvss.n3421 585
R2291 dvss.n3465 dvss.n3422 585
R2292 dvss.n3465 dvss.n3464 585
R2293 dvss.n3467 dvss.n3390 585
R2294 dvss.n3467 dvss.n3466 585
R2295 dvss.n3468 dvss.n3395 585
R2296 dvss.n3468 dvss.n3420 585
R2297 dvss.n3469 dvss.n3396 585
R2298 dvss.n3470 dvss.n3469 585
R2299 dvss.n3415 dvss.n3414 585
R2300 dvss.n3471 dvss.n3414 585
R2301 dvss.n3477 dvss.n3476 585
R2302 dvss.n3478 dvss.n3477 585
R2303 dvss.n3416 dvss.n3410 585
R2304 dvss.n3479 dvss.n3410 585
R2305 dvss.n3483 dvss.n3411 585
R2306 dvss.n3483 dvss.n3482 585
R2307 dvss.n3484 dvss.n3405 585
R2308 dvss.n3485 dvss.n3484 585
R2309 dvss.n3487 dvss.n3409 585
R2310 dvss.n3487 dvss.n3486 585
R2311 dvss.n3489 dvss.n3488 585
R2312 dvss.n3488 dvss.n121 585
R2313 dvss.n125 dvss.n122 585
R2314 dvss.n3649 dvss.n122 585
R2315 dvss.n1103 dvss.n1102 585
R2316 dvss.n624 dvss.n623 585
R2317 dvss.n1051 dvss.n1050 585
R2318 dvss.n630 dvss.n628 585
R2319 dvss.n1097 dvss.n1096 585
R2320 dvss.n1098 dvss.n1097 585
R2321 dvss.n1095 dvss.n629 585
R2322 dvss.n1061 dvss.n629 585
R2323 dvss.n1094 dvss.n1093 585
R2324 dvss.n1093 dvss.n1092 585
R2325 dvss.n635 dvss.n634 585
R2326 dvss.n1091 dvss.n635 585
R2327 dvss.n1089 dvss.n1088 585
R2328 dvss.n1090 dvss.n1089 585
R2329 dvss.n1087 dvss.n639 585
R2330 dvss.n646 dvss.n639 585
R2331 dvss.n1086 dvss.n1085 585
R2332 dvss.n1085 dvss.n1084 585
R2333 dvss.n644 dvss.n643 585
R2334 dvss.n672 dvss.n644 585
R2335 dvss.n671 dvss.n670 585
R2336 dvss.n675 dvss.n671 585
R2337 dvss.n678 dvss.n653 585
R2338 dvss.n678 dvss.n677 585
R2339 dvss.n679 dvss.n660 585
R2340 dvss.n680 dvss.n679 585
R2341 dvss.n668 dvss.n661 585
R2342 dvss.n681 dvss.n668 585
R2343 dvss.n685 dvss.n669 585
R2344 dvss.n685 dvss.n684 585
R2345 dvss.n686 dvss.n665 585
R2346 dvss.n687 dvss.n686 585
R2347 dvss.n569 dvss.n568 585
R2348 dvss.n688 dvss.n569 585
R2349 dvss.n1295 dvss.n1294 585
R2350 dvss.n1294 dvss.n1293 585
R2351 dvss.n562 dvss.n560 585
R2352 dvss.n560 dvss.n558 585
R2353 dvss.n1321 dvss.n1320 585
R2354 dvss.n1322 dvss.n1321 585
R2355 dvss.n1131 dvss.n1130 585
R2356 dvss.n1132 dvss.n1131 585
R2357 dvss.n603 dvss.n602 585
R2358 dvss.n1133 dvss.n603 585
R2359 dvss.n1136 dvss.n1135 585
R2360 dvss.n598 dvss.n597 585
R2361 dvss.n597 dvss.n596 585
R2362 dvss.n1146 dvss.n1145 585
R2363 dvss.n1147 dvss.n1146 585
R2364 dvss.n595 dvss.n594 585
R2365 dvss.n1152 dvss.n1151 585
R2366 dvss.n1151 dvss.n1150 585
R2367 dvss.n588 dvss.n587 585
R2368 dvss.n1149 dvss.n587 585
R2369 dvss.n1161 dvss.n1160 585
R2370 dvss.n1162 dvss.n1161 585
R2371 dvss.n586 dvss.n585 585
R2372 dvss.n1163 dvss.n586 585
R2373 dvss.n1167 dvss.n1166 585
R2374 dvss.n1166 dvss.n1165 585
R2375 dvss.n580 dvss.n579 585
R2376 dvss.n1164 dvss.n579 585
R2377 dvss.n1176 dvss.n1175 585
R2378 dvss.n1177 dvss.n1176 585
R2379 dvss.n578 dvss.n577 585
R2380 dvss.n1178 dvss.n578 585
R2381 dvss.n1181 dvss.n1180 585
R2382 dvss.n1180 dvss.n1179 585
R2383 dvss.n575 dvss.n573 585
R2384 dvss.n573 dvss.n571 585
R2385 dvss.n1289 dvss.n1288 585
R2386 dvss.n1290 dvss.n1289 585
R2387 dvss.n576 dvss.n574 585
R2388 dvss.n574 dvss.n572 585
R2389 dvss.n1284 dvss.n1184 585
R2390 dvss.n1283 dvss.n1185 585
R2391 dvss.n1212 dvss.n1186 585
R2392 dvss.n1279 dvss.n1187 585
R2393 dvss.n1278 dvss.n1188 585
R2394 dvss.n1217 dvss.n1188 585
R2395 dvss.n1219 dvss.n1189 585
R2396 dvss.n1219 dvss.n1218 585
R2397 dvss.n1220 dvss.n1192 585
R2398 dvss.n1270 dvss.n1193 585
R2399 dvss.n1222 dvss.n1193 585
R2400 dvss.n1269 dvss.n1194 585
R2401 dvss.n1223 dvss.n1194 585
R2402 dvss.n1211 dvss.n1195 585
R2403 dvss.n1261 dvss.n1199 585
R2404 dvss.n1227 dvss.n1199 585
R2405 dvss.n1260 dvss.n1200 585
R2406 dvss.n1228 dvss.n1200 585
R2407 dvss.n1229 dvss.n1201 585
R2408 dvss.n1230 dvss.n1229 585
R2409 dvss.n1253 dvss.n1203 585
R2410 dvss.n1231 dvss.n1203 585
R2411 dvss.n1252 dvss.n1204 585
R2412 dvss.n1232 dvss.n1204 585
R2413 dvss.n1234 dvss.n1205 585
R2414 dvss.n1234 dvss.n1233 585
R2415 dvss.n1235 dvss.n1209 585
R2416 dvss.n1236 dvss.n1235 585
R2417 dvss.n1243 dvss.n1210 585
R2418 dvss.n1237 dvss.n1210 585
R2419 dvss.n1242 dvss.n1239 585
R2420 dvss.n1239 dvss.n1238 585
R2421 dvss.n502 dvss.n501 585
R2422 dvss.n503 dvss.n502 585
R2423 dvss.n1586 dvss.n1585 585
R2424 dvss.n1585 dvss.n1584 585
R2425 dvss.n500 dvss.n499 585
R2426 dvss.n1583 dvss.n499 585
R2427 dvss.n1592 dvss.n1591 585
R2428 dvss.n498 dvss.n497 585
R2429 dvss.n1597 dvss.n1596 585
R2430 dvss.n496 dvss.n495 585
R2431 dvss.n1604 dvss.n1603 585
R2432 dvss.n1605 dvss.n1604 585
R2433 dvss.n493 dvss.n492 585
R2434 dvss.n1606 dvss.n493 585
R2435 dvss.n1609 dvss.n1608 585
R2436 dvss.n488 dvss.n487 585
R2437 dvss.n487 dvss.n486 585
R2438 dvss.n1619 dvss.n1618 585
R2439 dvss.n1620 dvss.n1619 585
R2440 dvss.n485 dvss.n484 585
R2441 dvss.n1625 dvss.n1624 585
R2442 dvss.n1624 dvss.n1623 585
R2443 dvss.n478 dvss.n477 585
R2444 dvss.n1622 dvss.n477 585
R2445 dvss.n1634 dvss.n1633 585
R2446 dvss.n1635 dvss.n1634 585
R2447 dvss.n476 dvss.n475 585
R2448 dvss.n1636 dvss.n476 585
R2449 dvss.n1640 dvss.n1639 585
R2450 dvss.n1639 dvss.n1638 585
R2451 dvss.n470 dvss.n469 585
R2452 dvss.n1637 dvss.n469 585
R2453 dvss.n1649 dvss.n1648 585
R2454 dvss.n1650 dvss.n1649 585
R2455 dvss.n468 dvss.n467 585
R2456 dvss.n1651 dvss.n468 585
R2457 dvss.n1654 dvss.n1653 585
R2458 dvss.n1653 dvss.n1652 585
R2459 dvss.n465 dvss.n463 585
R2460 dvss.n463 dvss.n461 585
R2461 dvss.n2879 dvss.n2878 585
R2462 dvss.n2880 dvss.n2879 585
R2463 dvss.n466 dvss.n464 585
R2464 dvss.n464 dvss.n462 585
R2465 dvss.n2874 dvss.n1657 585
R2466 dvss.n2873 dvss.n1658 585
R2467 dvss.n1792 dvss.n1659 585
R2468 dvss.n2869 dvss.n1660 585
R2469 dvss.n2868 dvss.n1661 585
R2470 dvss.n1797 dvss.n1661 585
R2471 dvss.n1799 dvss.n1662 585
R2472 dvss.n1799 dvss.n1798 585
R2473 dvss.n1800 dvss.n1665 585
R2474 dvss.n2860 dvss.n1666 585
R2475 dvss.n1802 dvss.n1666 585
R2476 dvss.n2859 dvss.n1667 585
R2477 dvss.n1803 dvss.n1667 585
R2478 dvss.n1791 dvss.n1668 585
R2479 dvss.n2851 dvss.n1672 585
R2480 dvss.n1807 dvss.n1672 585
R2481 dvss.n2850 dvss.n1673 585
R2482 dvss.n1808 dvss.n1673 585
R2483 dvss.n1809 dvss.n1674 585
R2484 dvss.n1810 dvss.n1809 585
R2485 dvss.n2843 dvss.n1676 585
R2486 dvss.n1811 dvss.n1676 585
R2487 dvss.n2842 dvss.n1677 585
R2488 dvss.n1812 dvss.n1677 585
R2489 dvss.n1814 dvss.n1678 585
R2490 dvss.n1814 dvss.n1813 585
R2491 dvss.n1815 dvss.n1682 585
R2492 dvss.n1816 dvss.n1815 585
R2493 dvss.n2833 dvss.n1683 585
R2494 dvss.n1817 dvss.n1683 585
R2495 dvss.n2832 dvss.n1684 585
R2496 dvss.n1818 dvss.n1684 585
R2497 dvss.n1819 dvss.n1685 585
R2498 dvss.n1820 dvss.n1819 585
R2499 dvss.n2828 dvss.n1686 585
R2500 dvss.n1822 dvss.n1686 585
R2501 dvss.n2827 dvss.n1687 585
R2502 dvss.n1823 dvss.n1687 585
R2503 dvss.n1788 dvss.n1688 585
R2504 dvss.n2823 dvss.n1689 585
R2505 dvss.n2822 dvss.n1690 585
R2506 dvss.n1786 dvss.n1691 585
R2507 dvss.n2818 dvss.n1692 585
R2508 dvss.n1825 dvss.n1692 585
R2509 dvss.n2817 dvss.n1693 585
R2510 dvss.n1826 dvss.n1693 585
R2511 dvss.n1827 dvss.n1694 585
R2512 dvss.n2810 dvss.n1697 585
R2513 dvss.n1829 dvss.n1697 585
R2514 dvss.n2809 dvss.n1698 585
R2515 dvss.n1830 dvss.n1698 585
R2516 dvss.n1785 dvss.n1699 585
R2517 dvss.n2801 dvss.n1703 585
R2518 dvss.n1832 dvss.n1703 585
R2519 dvss.n2800 dvss.n1704 585
R2520 dvss.n1833 dvss.n1704 585
R2521 dvss.n1834 dvss.n1705 585
R2522 dvss.n1835 dvss.n1834 585
R2523 dvss.n2793 dvss.n1707 585
R2524 dvss.n1836 dvss.n1707 585
R2525 dvss.n2792 dvss.n1708 585
R2526 dvss.n1837 dvss.n1708 585
R2527 dvss.n1839 dvss.n1709 585
R2528 dvss.n1839 dvss.n1838 585
R2529 dvss.n1840 dvss.n1713 585
R2530 dvss.n1841 dvss.n1840 585
R2531 dvss.n2783 dvss.n1714 585
R2532 dvss.n1842 dvss.n1714 585
R2533 dvss.n2782 dvss.n1715 585
R2534 dvss.n1843 dvss.n1715 585
R2535 dvss.n1844 dvss.n1716 585
R2536 dvss.n1845 dvss.n1844 585
R2537 dvss.n2778 dvss.n1717 585
R2538 dvss.n1847 dvss.n1717 585
R2539 dvss.n2777 dvss.n1718 585
R2540 dvss.n1848 dvss.n1718 585
R2541 dvss.n1782 dvss.n1719 585
R2542 dvss.n2773 dvss.n1720 585
R2543 dvss.n2772 dvss.n1721 585
R2544 dvss.n1780 dvss.n1722 585
R2545 dvss.n2768 dvss.n1723 585
R2546 dvss.n1850 dvss.n1723 585
R2547 dvss.n2767 dvss.n1724 585
R2548 dvss.n1851 dvss.n1724 585
R2549 dvss.n1852 dvss.n1725 585
R2550 dvss.n2760 dvss.n1728 585
R2551 dvss.n1854 dvss.n1728 585
R2552 dvss.n2759 dvss.n1729 585
R2553 dvss.n1855 dvss.n1729 585
R2554 dvss.n1779 dvss.n1730 585
R2555 dvss.n2751 dvss.n1734 585
R2556 dvss.n1857 dvss.n1734 585
R2557 dvss.n2750 dvss.n1735 585
R2558 dvss.n1858 dvss.n1735 585
R2559 dvss.n1859 dvss.n1736 585
R2560 dvss.n1860 dvss.n1859 585
R2561 dvss.n2743 dvss.n1738 585
R2562 dvss.n1861 dvss.n1738 585
R2563 dvss.n2742 dvss.n1739 585
R2564 dvss.n1862 dvss.n1739 585
R2565 dvss.n1864 dvss.n1740 585
R2566 dvss.n1864 dvss.n1863 585
R2567 dvss.n1865 dvss.n1744 585
R2568 dvss.n1866 dvss.n1865 585
R2569 dvss.n2733 dvss.n1745 585
R2570 dvss.n1867 dvss.n1745 585
R2571 dvss.n2732 dvss.n1746 585
R2572 dvss.n1868 dvss.n1746 585
R2573 dvss.n1869 dvss.n1747 585
R2574 dvss.n1870 dvss.n1869 585
R2575 dvss.n2728 dvss.n1748 585
R2576 dvss.n1872 dvss.n1748 585
R2577 dvss.n2727 dvss.n1749 585
R2578 dvss.n1873 dvss.n1749 585
R2579 dvss.n1876 dvss.n1750 585
R2580 dvss.n2723 dvss.n1751 585
R2581 dvss.n2722 dvss.n1752 585
R2582 dvss.n1874 dvss.n1753 585
R2583 dvss.n2718 dvss.n1754 585
R2584 dvss.n1880 dvss.n1754 585
R2585 dvss.n2717 dvss.n1755 585
R2586 dvss.n1881 dvss.n1755 585
R2587 dvss.n1882 dvss.n1756 585
R2588 dvss.n2710 dvss.n1759 585
R2589 dvss.n1884 dvss.n1759 585
R2590 dvss.n2709 dvss.n1760 585
R2591 dvss.n1885 dvss.n1760 585
R2592 dvss.n1778 dvss.n1761 585
R2593 dvss.n2701 dvss.n1765 585
R2594 dvss.n2672 dvss.n1765 585
R2595 dvss.n2700 dvss.n1766 585
R2596 dvss.n2673 dvss.n1766 585
R2597 dvss.n2674 dvss.n1767 585
R2598 dvss.n2675 dvss.n2674 585
R2599 dvss.n2693 dvss.n1769 585
R2600 dvss.n2676 dvss.n1769 585
R2601 dvss.n2692 dvss.n1770 585
R2602 dvss.n2677 dvss.n1770 585
R2603 dvss.n2678 dvss.n1771 585
R2604 dvss.n2679 dvss.n2678 585
R2605 dvss.n1777 dvss.n1776 585
R2606 dvss.n2680 dvss.n1777 585
R2607 dvss.n2683 dvss.n2682 585
R2608 dvss.n2682 dvss.n2681 585
R2609 dvss.n169 dvss.n168 585
R2610 dvss.n170 dvss.n169 585
R2611 dvss.n3551 dvss.n3550 585
R2612 dvss.n3550 dvss.n3549 585
R2613 dvss.n166 dvss.n164 585
R2614 dvss.n164 dvss.n163 585
R2615 dvss.n3569 dvss.n3568 585
R2616 dvss.n3570 dvss.n3569 585
R2617 dvss.n167 dvss.n165 585
R2618 dvss.n3564 dvss.n3555 585
R2619 dvss.n3563 dvss.n3556 585
R2620 dvss.n3559 dvss.n3558 585
R2621 dvss.n161 dvss.n160 585
R2622 dvss.n3572 dvss.n161 585
R2623 dvss.n3576 dvss.n3575 585
R2624 dvss.n3575 dvss.n3574 585
R2625 dvss.n157 dvss.n156 585
R2626 dvss.n3588 dvss.n3587 585
R2627 dvss.n3589 dvss.n3588 585
R2628 dvss.n155 dvss.n154 585
R2629 dvss.n3590 dvss.n155 585
R2630 dvss.n3593 dvss.n3592 585
R2631 dvss.n149 dvss.n148 585
R2632 dvss.n148 dvss.n147 585
R2633 dvss.n3603 dvss.n3602 585
R2634 dvss.n3604 dvss.n3603 585
R2635 dvss.n145 dvss.n144 585
R2636 dvss.n3605 dvss.n145 585
R2637 dvss.n3608 dvss.n3607 585
R2638 dvss.n3607 dvss.n3606 585
R2639 dvss.n143 dvss.n142 585
R2640 dvss.n142 dvss.n141 585
R2641 dvss.n3621 dvss.n3620 585
R2642 dvss.n3622 dvss.n3621 585
R2643 dvss.n140 dvss.n139 585
R2644 dvss.n3623 dvss.n140 585
R2645 dvss.n3626 dvss.n3625 585
R2646 dvss.n3625 dvss.n3624 585
R2647 dvss.n137 dvss.n136 585
R2648 dvss.n136 dvss.n135 585
R2649 dvss.n3634 dvss.n3633 585
R2650 dvss.n3635 dvss.n3634 585
R2651 dvss.n138 dvss.n132 585
R2652 dvss.n3637 dvss.n132 585
R2653 dvss.n3639 dvss.n133 585
R2654 dvss.n3639 dvss.n3638 585
R2655 dvss.n3640 dvss.n131 585
R2656 dvss.n1119 dvss.n1118 585
R2657 dvss.n608 dvss.n607 585
R2658 dvss.n1124 dvss.n1123 585
R2659 dvss.n606 dvss.n605 585
R2660 dvss.n852 dvss.n851 585
R2661 dvss.n851 dvss.n765 585
R2662 dvss.n850 dvss.n771 585
R2663 dvss.n850 dvss.n849 585
R2664 dvss.n775 dvss.n772 585
R2665 dvss.n846 dvss.n845 585
R2666 dvss.n847 dvss.n846 585
R2667 dvss.n844 dvss.n774 585
R2668 dvss.n774 dvss.n773 585
R2669 dvss.n843 dvss.n842 585
R2670 dvss.n780 dvss.n779 585
R2671 dvss.n840 dvss.n780 585
R2672 dvss.n838 dvss.n837 585
R2673 dvss.n839 dvss.n838 585
R2674 dvss.n836 dvss.n781 585
R2675 dvss.n806 dvss.n781 585
R2676 dvss.n835 dvss.n834 585
R2677 dvss.n834 dvss.n833 585
R2678 dvss.n805 dvss.n804 585
R2679 dvss.n832 dvss.n805 585
R2680 dvss.n830 dvss.n829 585
R2681 dvss.n831 dvss.n830 585
R2682 dvss.n828 dvss.n807 585
R2683 dvss.n823 dvss.n807 585
R2684 dvss.n827 dvss.n826 585
R2685 dvss.n826 dvss.n825 585
R2686 dvss.n822 dvss.n821 585
R2687 dvss.n824 dvss.n822 585
R2688 dvss.n612 dvss.n611 585
R2689 dvss.n613 dvss.n612 585
R2690 dvss.n1113 dvss.n1112 585
R2691 dvss.n1112 dvss.n1111 585
R2692 dvss.n610 dvss.n609 585
R2693 dvss.n1110 dvss.n609 585
R2694 dvss.n988 dvss.n985 585
R2695 dvss.n988 dvss.n987 585
R2696 dvss.n739 dvss.n736 585
R2697 dvss.n1003 dvss.n739 585
R2698 dvss.n1007 dvss.n1006 585
R2699 dvss.n1006 dvss.n1005 585
R2700 dvss.n1008 dvss.n731 585
R2701 dvss.n733 dvss.n731 585
R2702 dvss.n1021 dvss.n732 585
R2703 dvss.n1021 dvss.n1020 585
R2704 dvss.n1022 dvss.n724 585
R2705 dvss.n1023 dvss.n1022 585
R2706 dvss.n730 dvss.n729 585
R2707 dvss.n1024 dvss.n730 585
R2708 dvss.n1028 dvss.n1027 585
R2709 dvss.n1027 dvss.n1026 585
R2710 dvss.n619 dvss.n617 585
R2711 dvss.n617 dvss.n614 585
R2712 dvss.n1106 dvss.n1105 585
R2713 dvss.n1107 dvss.n1106 585
R2714 dvss.n1104 dvss.n618 585
R2715 dvss.n618 dvss.n616 585
R2716 dvss.n961 dvss.n960 585
R2717 dvss.n960 dvss.n959 585
R2718 dvss.n962 dvss.n759 585
R2719 dvss.n857 dvss.n759 585
R2720 dvss.n969 dvss.n758 585
R2721 dvss.n969 dvss.n968 585
R2722 dvss.n971 dvss.n970 585
R2723 dvss.n970 dvss.n751 585
R2724 dvss.n754 dvss.n749 585
R2725 dvss.n981 dvss.n749 585
R2726 dvss.n983 dvss.n750 585
R2727 dvss.n983 dvss.n982 585
R2728 dvss.n989 dvss.n745 585
R2729 dvss.n990 dvss.n989 585
R2730 dvss.n958 dvss.n957 585
R2731 dvss.n959 dvss.n958 585
R2732 dvss.n761 dvss.n760 585
R2733 dvss.n857 dvss.n760 585
R2734 dvss.n967 dvss.n966 585
R2735 dvss.n968 dvss.n967 585
R2736 dvss.n753 dvss.n752 585
R2737 dvss.n752 dvss.n751 585
R2738 dvss.n980 dvss.n979 585
R2739 dvss.n981 dvss.n980 585
R2740 dvss.n747 dvss.n746 585
R2741 dvss.n982 dvss.n747 585
R2742 dvss.n992 dvss.n991 585
R2743 dvss.n991 dvss.n990 585
R2744 dvss.n741 dvss.n740 585
R2745 dvss.n987 dvss.n740 585
R2746 dvss.n1002 dvss.n1001 585
R2747 dvss.n1003 dvss.n1002 585
R2748 dvss.n735 dvss.n734 585
R2749 dvss.n1005 dvss.n734 585
R2750 dvss.n1018 dvss.n1017 585
R2751 dvss.n1018 dvss.n733 585
R2752 dvss.n1019 dvss.n726 585
R2753 dvss.n1020 dvss.n1019 585
R2754 dvss.n1032 dvss.n727 585
R2755 dvss.n1023 dvss.n727 585
R2756 dvss.n1031 dvss.n728 585
R2757 dvss.n1024 dvss.n728 585
R2758 dvss.n1025 dvss.n718 585
R2759 dvss.n1026 dvss.n1025 585
R2760 dvss.n1041 dvss.n719 585
R2761 dvss.n719 dvss.n614 585
R2762 dvss.n1042 dvss.n615 585
R2763 dvss.n1107 dvss.n615 585
R2764 dvss.n1044 dvss.n1043 585
R2765 dvss.n1044 dvss.n616 585
R2766 dvss.n1045 dvss.n714 585
R2767 dvss.n1048 dvss.n1047 585
R2768 dvss.n715 dvss.n712 585
R2769 dvss.n1059 dvss.n713 585
R2770 dvss.n1060 dvss.n627 585
R2771 dvss.n1098 dvss.n627 585
R2772 dvss.n1063 dvss.n1062 585
R2773 dvss.n1062 dvss.n1061 585
R2774 dvss.n1064 dvss.n636 585
R2775 dvss.n1092 dvss.n636 585
R2776 dvss.n1066 dvss.n637 585
R2777 dvss.n1091 dvss.n637 585
R2778 dvss.n1065 dvss.n638 585
R2779 dvss.n1090 dvss.n638 585
R2780 dvss.n649 dvss.n647 585
R2781 dvss.n647 dvss.n646 585
R2782 dvss.n1083 dvss.n1082 585
R2783 dvss.n1084 dvss.n1083 585
R2784 dvss.n1081 dvss.n648 585
R2785 dvss.n672 dvss.n648 585
R2786 dvss.n674 dvss.n650 585
R2787 dvss.n675 dvss.n674 585
R2788 dvss.n706 dvss.n654 585
R2789 dvss.n677 dvss.n654 585
R2790 dvss.n705 dvss.n655 585
R2791 dvss.n680 dvss.n655 585
R2792 dvss.n682 dvss.n656 585
R2793 dvss.n682 dvss.n681 585
R2794 dvss.n683 dvss.n666 585
R2795 dvss.n684 dvss.n683 585
R2796 dvss.n692 dvss.n667 585
R2797 dvss.n687 dvss.n667 585
R2798 dvss.n691 dvss.n689 585
R2799 dvss.n689 dvss.n688 585
R2800 dvss.n570 dvss.n565 585
R2801 dvss.n1293 dvss.n570 585
R2802 dvss.n1301 dvss.n566 585
R2803 dvss.n566 dvss.n558 585
R2804 dvss.n1302 dvss.n559 585
R2805 dvss.n1322 dvss.n559 585
R2806 dvss.n1317 dvss.n1303 585
R2807 dvss.n1316 dvss.n1308 585
R2808 dvss.n1304 dvss.n554 585
R2809 dvss.n1327 dvss.n555 585
R2810 dvss.n1326 dvss.n1325 585
R2811 dvss.n1325 dvss.n1324 585
R2812 dvss.n549 dvss.n548 585
R2813 dvss.n1337 dvss.n549 585
R2814 dvss.n1340 dvss.n1339 585
R2815 dvss.n1339 dvss.n1338 585
R2816 dvss.n543 dvss.n542 585
R2817 dvss.n544 dvss.n543 585
R2818 dvss.n1353 dvss.n1352 585
R2819 dvss.n1352 dvss.n1351 585
R2820 dvss.n538 dvss.n537 585
R2821 dvss.n545 dvss.n537 585
R2822 dvss.n1368 dvss.n1367 585
R2823 dvss.n1369 dvss.n1368 585
R2824 dvss.n534 dvss.n533 585
R2825 dvss.n1372 dvss.n534 585
R2826 dvss.n1377 dvss.n1376 585
R2827 dvss.n1376 dvss.n1375 585
R2828 dvss.n529 dvss.n528 585
R2829 dvss.n1225 dvss.n528 585
R2830 dvss.n1395 dvss.n1394 585
R2831 dvss.n1395 dvss.n527 585
R2832 dvss.n1396 dvss.n520 585
R2833 dvss.n1397 dvss.n1396 585
R2834 dvss.n1409 dvss.n521 585
R2835 dvss.n1400 dvss.n521 585
R2836 dvss.n1408 dvss.n522 585
R2837 dvss.n1401 dvss.n522 585
R2838 dvss.n1402 dvss.n512 585
R2839 dvss.n1403 dvss.n1402 585
R2840 dvss.n1417 dvss.n513 585
R2841 dvss.n513 dvss.n504 585
R2842 dvss.n1576 dvss.n505 585
R2843 dvss.n1580 dvss.n505 585
R2844 dvss.n1575 dvss.n1418 585
R2845 dvss.n1418 dvss.n506 585
R2846 dvss.n1478 dvss.n1419 585
R2847 dvss.n1571 dvss.n1422 585
R2848 dvss.n1570 dvss.n1423 585
R2849 dvss.n1482 dvss.n1424 585
R2850 dvss.n1483 dvss.n1431 585
R2851 dvss.n1493 dvss.n1483 585
R2852 dvss.n1563 dvss.n1432 585
R2853 dvss.n1494 dvss.n1432 585
R2854 dvss.n1562 dvss.n1433 585
R2855 dvss.n1495 dvss.n1433 585
R2856 dvss.n1473 dvss.n1434 585
R2857 dvss.n1473 dvss.n1472 585
R2858 dvss.n1474 dvss.n1442 585
R2859 dvss.n1503 dvss.n1474 585
R2860 dvss.n1554 dvss.n1443 585
R2861 dvss.n1504 dvss.n1443 585
R2862 dvss.n1553 dvss.n1444 585
R2863 dvss.n1506 dvss.n1444 585
R2864 dvss.n1510 dvss.n1445 585
R2865 dvss.n1510 dvss.n1509 585
R2866 dvss.n1511 dvss.n1451 585
R2867 dvss.n1512 dvss.n1511 585
R2868 dvss.n1543 dvss.n1452 585
R2869 dvss.n1514 dvss.n1452 585
R2870 dvss.n1542 dvss.n1453 585
R2871 dvss.n1517 dvss.n1453 585
R2872 dvss.n1519 dvss.n1454 585
R2873 dvss.n1519 dvss.n1518 585
R2874 dvss.n1520 dvss.n1464 585
R2875 dvss.n1521 dvss.n1520 585
R2876 dvss.n1529 dvss.n1465 585
R2877 dvss.n1524 dvss.n1465 585
R2878 dvss.n1528 dvss.n1526 585
R2879 dvss.n1526 dvss.n1525 585
R2880 dvss.n460 dvss.n455 585
R2881 dvss.n2883 dvss.n460 585
R2882 dvss.n2891 dvss.n456 585
R2883 dvss.n456 dvss.n449 585
R2884 dvss.n2910 dvss.n450 585
R2885 dvss.n2914 dvss.n450 585
R2886 dvss.n2909 dvss.n2892 585
R2887 dvss.n2898 dvss.n2897 585
R2888 dvss.n2893 dvss.n445 585
R2889 dvss.n2919 dvss.n446 585
R2890 dvss.n2918 dvss.n2917 585
R2891 dvss.n2917 dvss.n2916 585
R2892 dvss.n440 dvss.n439 585
R2893 dvss.n2929 dvss.n440 585
R2894 dvss.n2932 dvss.n2931 585
R2895 dvss.n2931 dvss.n2930 585
R2896 dvss.n434 dvss.n433 585
R2897 dvss.n435 dvss.n434 585
R2898 dvss.n2945 dvss.n2944 585
R2899 dvss.n2944 dvss.n2943 585
R2900 dvss.n429 dvss.n428 585
R2901 dvss.n436 dvss.n428 585
R2902 dvss.n2960 dvss.n2959 585
R2903 dvss.n2961 dvss.n2960 585
R2904 dvss.n425 dvss.n424 585
R2905 dvss.n2964 dvss.n425 585
R2906 dvss.n2969 dvss.n2968 585
R2907 dvss.n2968 dvss.n2967 585
R2908 dvss.n420 dvss.n419 585
R2909 dvss.n1805 dvss.n419 585
R2910 dvss.n2987 dvss.n2986 585
R2911 dvss.n2987 dvss.n418 585
R2912 dvss.n2988 dvss.n411 585
R2913 dvss.n2989 dvss.n2988 585
R2914 dvss.n3002 dvss.n412 585
R2915 dvss.n2992 dvss.n412 585
R2916 dvss.n3001 dvss.n413 585
R2917 dvss.n2993 dvss.n413 585
R2918 dvss.n2994 dvss.n403 585
R2919 dvss.n2996 dvss.n2994 585
R2920 dvss.n3010 dvss.n404 585
R2921 dvss.n2995 dvss.n404 585
R2922 dvss.n3011 dvss.n397 585
R2923 dvss.n3015 dvss.n397 585
R2924 dvss.n3017 dvss.n396 585
R2925 dvss.n3017 dvss.n3016 585
R2926 dvss.n3030 dvss.n3018 585
R2927 dvss.n3029 dvss.n3019 585
R2928 dvss.n3026 dvss.n3025 585
R2929 dvss.n3020 dvss.n386 585
R2930 dvss.n3046 dvss.n387 585
R2931 dvss.n390 dvss.n387 585
R2932 dvss.n3047 dvss.n380 585
R2933 dvss.n3051 dvss.n380 585
R2934 dvss.n3053 dvss.n381 585
R2935 dvss.n3053 dvss.n3052 585
R2936 dvss.n3054 dvss.n374 585
R2937 dvss.n3056 dvss.n3054 585
R2938 dvss.n3072 dvss.n375 585
R2939 dvss.n3055 dvss.n375 585
R2940 dvss.n3073 dvss.n371 585
R2941 dvss.n3077 dvss.n371 585
R2942 dvss.n370 dvss.n364 585
R2943 dvss.n370 dvss.n369 585
R2944 dvss.n3084 dvss.n365 585
R2945 dvss.n3080 dvss.n365 585
R2946 dvss.n3085 dvss.n359 585
R2947 dvss.n368 dvss.n359 585
R2948 dvss.n3095 dvss.n358 585
R2949 dvss.n3095 dvss.n3094 585
R2950 dvss.n3097 dvss.n3096 585
R2951 dvss.n3096 dvss.n354 585
R2952 dvss.n355 dvss.n348 585
R2953 dvss.n3108 dvss.n355 585
R2954 dvss.n3119 dvss.n349 585
R2955 dvss.n3109 dvss.n349 585
R2956 dvss.n3118 dvss.n350 585
R2957 dvss.n3113 dvss.n350 585
R2958 dvss.n3110 dvss.n351 585
R2959 dvss.n3112 dvss.n3110 585
R2960 dvss.n338 dvss.n337 585
R2961 dvss.n3111 dvss.n337 585
R2962 dvss.n3132 dvss.n3131 585
R2963 dvss.n3133 dvss.n3132 585
R2964 dvss.n326 dvss.n325 585
R2965 dvss.n3134 dvss.n325 585
R2966 dvss.n3146 dvss.n3145 585
R2967 dvss.n327 dvss.n324 585
R2968 dvss.n322 dvss.n321 585
R2969 dvss.n3152 dvss.n3150 585
R2970 dvss.n3151 dvss.n315 585
R2971 dvss.n332 dvss.n315 585
R2972 dvss.n3169 dvss.n316 585
R2973 dvss.n3169 dvss.n3168 585
R2974 dvss.n3170 dvss.n311 585
R2975 dvss.n3171 dvss.n3170 585
R2976 dvss.n3177 dvss.n312 585
R2977 dvss.n3173 dvss.n312 585
R2978 dvss.n3178 dvss.n305 585
R2979 dvss.n3172 dvss.n305 585
R2980 dvss.n3191 dvss.n306 585
R2981 dvss.n3191 dvss.n3190 585
R2982 dvss.n3192 dvss.n300 585
R2983 dvss.n3193 dvss.n3192 585
R2984 dvss.n3200 dvss.n301 585
R2985 dvss.n3196 dvss.n301 585
R2986 dvss.n3201 dvss.n295 585
R2987 dvss.n304 dvss.n295 585
R2988 dvss.n3211 dvss.n294 585
R2989 dvss.n3211 dvss.n3210 585
R2990 dvss.n3213 dvss.n3212 585
R2991 dvss.n3212 dvss.n290 585
R2992 dvss.n291 dvss.n284 585
R2993 dvss.n3224 dvss.n291 585
R2994 dvss.n3235 dvss.n285 585
R2995 dvss.n3225 dvss.n285 585
R2996 dvss.n3234 dvss.n286 585
R2997 dvss.n3229 dvss.n286 585
R2998 dvss.n3226 dvss.n287 585
R2999 dvss.n3228 dvss.n3226 585
R3000 dvss.n274 dvss.n273 585
R3001 dvss.n3227 dvss.n273 585
R3002 dvss.n3248 dvss.n3247 585
R3003 dvss.n3249 dvss.n3248 585
R3004 dvss.n262 dvss.n261 585
R3005 dvss.n3250 dvss.n261 585
R3006 dvss.n3262 dvss.n3261 585
R3007 dvss.n263 dvss.n260 585
R3008 dvss.n258 dvss.n257 585
R3009 dvss.n3267 dvss.n3266 585
R3010 dvss.n254 dvss.n253 585
R3011 dvss.n268 dvss.n253 585
R3012 dvss.n3285 dvss.n3284 585
R3013 dvss.n3286 dvss.n3285 585
R3014 dvss.n248 dvss.n247 585
R3015 dvss.n3287 dvss.n248 585
R3016 dvss.n3292 dvss.n3291 585
R3017 dvss.n3291 dvss.n3290 585
R3018 dvss.n249 dvss.n243 585
R3019 dvss.n250 dvss.n249 585
R3020 dvss.n3305 dvss.n239 585
R3021 dvss.n3309 dvss.n239 585
R3022 dvss.n3304 dvss.n244 585
R3023 dvss.n244 dvss.n238 585
R3024 dvss.n235 dvss.n234 585
R3025 dvss.n3312 dvss.n235 585
R3026 dvss.n3317 dvss.n3316 585
R3027 dvss.n3316 dvss.n3315 585
R3028 dvss.n230 dvss.n229 585
R3029 dvss.n1887 dvss.n229 585
R3030 dvss.n3335 dvss.n3334 585
R3031 dvss.n3335 dvss.n228 585
R3032 dvss.n3336 dvss.n221 585
R3033 dvss.n3337 dvss.n3336 585
R3034 dvss.n3349 dvss.n222 585
R3035 dvss.n3340 dvss.n222 585
R3036 dvss.n3348 dvss.n223 585
R3037 dvss.n3341 dvss.n223 585
R3038 dvss.n3342 dvss.n213 585
R3039 dvss.n3343 dvss.n3342 585
R3040 dvss.n3357 dvss.n214 585
R3041 dvss.n214 dvss.n205 585
R3042 dvss.n3542 dvss.n206 585
R3043 dvss.n3546 dvss.n206 585
R3044 dvss.n3541 dvss.n3358 585
R3045 dvss.n3358 dvss.n207 585
R3046 dvss.n3440 dvss.n3359 585
R3047 dvss.n3537 dvss.n3362 585
R3048 dvss.n3536 dvss.n3363 585
R3049 dvss.n3444 dvss.n3364 585
R3050 dvss.n3445 dvss.n3371 585
R3051 dvss.n3446 dvss.n3445 585
R3052 dvss.n3529 dvss.n3372 585
R3053 dvss.n3447 dvss.n3372 585
R3054 dvss.n3528 dvss.n3373 585
R3055 dvss.n3450 dvss.n3373 585
R3056 dvss.n3452 dvss.n3374 585
R3057 dvss.n3452 dvss.n3451 585
R3058 dvss.n3453 dvss.n3382 585
R3059 dvss.n3454 dvss.n3453 585
R3060 dvss.n3520 dvss.n3383 585
R3061 dvss.n3458 dvss.n3383 585
R3062 dvss.n3519 dvss.n3384 585
R3063 dvss.n3423 dvss.n3384 585
R3064 dvss.n3462 dvss.n3385 585
R3065 dvss.n3462 dvss.n3461 585
R3066 dvss.n3463 dvss.n3391 585
R3067 dvss.n3464 dvss.n3463 585
R3068 dvss.n3509 dvss.n3392 585
R3069 dvss.n3466 dvss.n3392 585
R3070 dvss.n3508 dvss.n3393 585
R3071 dvss.n3420 dvss.n3393 585
R3072 dvss.n3419 dvss.n3394 585
R3073 dvss.n3470 dvss.n3419 585
R3074 dvss.n3473 dvss.n3472 585
R3075 dvss.n3472 dvss.n3471 585
R3076 dvss.n3474 dvss.n3412 585
R3077 dvss.n3478 dvss.n3412 585
R3078 dvss.n3480 dvss.n3413 585
R3079 dvss.n3480 dvss.n3479 585
R3080 dvss.n3481 dvss.n3406 585
R3081 dvss.n3482 dvss.n3481 585
R3082 dvss.n3493 dvss.n3407 585
R3083 dvss.n3485 dvss.n3407 585
R3084 dvss.n3492 dvss.n3408 585
R3085 dvss.n3486 dvss.n3408 585
R3086 dvss.n124 dvss.n123 585
R3087 dvss.n123 dvss.n121 585
R3088 dvss.n3648 dvss.n3647 585
R3089 dvss.n3649 dvss.n3648 585
R3090 dvss.n956 dvss.n858 585
R3091 dvss.n945 dvss.n862 585
R3092 dvss.n948 dvss.n947 585
R3093 dvss.n764 dvss.n762 585
R3094 dvss.n863 dvss.n764 585
R3095 dvss.n853 dvss.n766 585
R3096 dvss.n899 dvss.n898 585
R3097 dvss.n900 dvss.n899 585
R3098 dvss.n897 dvss.n877 585
R3099 dvss.n877 dvss.n876 585
R3100 dvss.n896 dvss.n895 585
R3101 dvss.n895 dvss.n894 585
R3102 dvss.n881 dvss.n880 585
R3103 dvss.n893 dvss.n881 585
R3104 dvss.n891 dvss.n890 585
R3105 dvss.n892 dvss.n891 585
R3106 dvss.n889 dvss.n883 585
R3107 dvss.n883 dvss.n882 585
R3108 dvss.n874 dvss.n873 585
R3109 dvss.n875 dvss.n874 585
R3110 dvss.n908 dvss.n907 585
R3111 dvss.n907 dvss.n906 585
R3112 dvss.n872 dvss.n871 585
R3113 dvss.n904 dvss.n871 585
R3114 dvss.n921 dvss.n920 585
R3115 dvss.n922 dvss.n921 585
R3116 dvss.n870 dvss.n869 585
R3117 dvss.n923 dvss.n870 585
R3118 dvss.n927 dvss.n926 585
R3119 dvss.n926 dvss.n925 585
R3120 dvss.n867 dvss.n866 585
R3121 dvss.n924 dvss.n866 585
R3122 dvss.n940 dvss.n939 585
R3123 dvss.n941 dvss.n940 585
R3124 dvss.n938 dvss.n864 585
R3125 dvss.n942 dvss.n864 585
R3126 dvss.n944 dvss.n865 585
R3127 dvss.n944 dvss.n943 585
R3128 dvss.n2665 dvss.n2664 585
R3129 dvss.n2666 dvss.n2665 585
R3130 dvss.n1966 dvss.n1965 585
R3131 dvss.n2661 dvss.n1967 585
R3132 dvss.n2660 dvss.n1968 585
R3133 dvss.n1970 dvss.n1969 585
R3134 dvss.n2655 dvss.n1971 585
R3135 dvss.n2654 dvss.n1972 585
R3136 dvss.n1974 dvss.n1973 585
R3137 dvss.n2650 dvss.n1975 585
R3138 dvss.n2649 dvss.n1976 585
R3139 dvss.n1981 dvss.n1977 585
R3140 dvss.n2642 dvss.n1982 585
R3141 dvss.n2641 dvss.n1983 585
R3142 dvss.n1985 dvss.n1984 585
R3143 dvss.n1991 dvss.n1990 585
R3144 dvss.n2634 dvss.n1992 585
R3145 dvss.n2633 dvss.n1993 585
R3146 dvss.n2630 dvss.n1994 585
R3147 dvss.n2629 dvss.n1995 585
R3148 dvss.n1997 dvss.n1996 585
R3149 dvss.n2623 dvss.n2001 585
R3150 dvss.n2622 dvss.n2002 585
R3151 dvss.n2004 dvss.n2003 585
R3152 dvss.n2618 dvss.n2005 585
R3153 dvss.n2617 dvss.n2006 585
R3154 dvss.n2008 dvss.n2007 585
R3155 dvss.n2613 dvss.n2009 585
R3156 dvss.n2612 dvss.n2010 585
R3157 dvss.n2014 dvss.n2011 585
R3158 dvss.n2605 dvss.n2015 585
R3159 dvss.n2604 dvss.n2016 585
R3160 dvss.n2018 dvss.n2017 585
R3161 dvss.n2597 dvss.n2020 585
R3162 dvss.n2596 dvss.n2021 585
R3163 dvss.n2023 dvss.n2022 585
R3164 dvss.n2589 dvss.n2024 585
R3165 dvss.n2588 dvss.n2025 585
R3166 dvss.n2027 dvss.n2026 585
R3167 dvss.n2584 dvss.n2028 585
R3168 dvss.n2583 dvss.n2029 585
R3169 dvss.n2034 dvss.n2030 585
R3170 dvss.n2036 dvss.n2035 585
R3171 dvss.n2576 dvss.n2037 585
R3172 dvss.n2575 dvss.n2038 585
R3173 dvss.n2040 dvss.n2039 585
R3174 dvss.n2571 dvss.n2041 585
R3175 dvss.n2570 dvss.n2042 585
R3176 dvss.n2044 dvss.n2043 585
R3177 dvss.n2566 dvss.n2045 585
R3178 dvss.n2565 dvss.n2046 585
R3179 dvss.n2050 dvss.n2047 585
R3180 dvss.n2558 dvss.n2051 585
R3181 dvss.n2557 dvss.n2052 585
R3182 dvss.n2054 dvss.n2053 585
R3183 dvss.n2550 dvss.n2056 585
R3184 dvss.n2549 dvss.n2057 585
R3185 dvss.n2059 dvss.n2058 585
R3186 dvss.n2542 dvss.n2060 585
R3187 dvss.n2541 dvss.n2061 585
R3188 dvss.n2063 dvss.n2062 585
R3189 dvss.n2537 dvss.n2064 585
R3190 dvss.n2536 dvss.n2065 585
R3191 dvss.n2070 dvss.n2066 585
R3192 dvss.n2072 dvss.n2071 585
R3193 dvss.n2529 dvss.n2073 585
R3194 dvss.n2528 dvss.n2074 585
R3195 dvss.n2076 dvss.n2075 585
R3196 dvss.n2524 dvss.n2077 585
R3197 dvss.n2523 dvss.n2078 585
R3198 dvss.n2080 dvss.n2079 585
R3199 dvss.n2519 dvss.n2081 585
R3200 dvss.n2518 dvss.n2082 585
R3201 dvss.n2086 dvss.n2083 585
R3202 dvss.n2511 dvss.n2087 585
R3203 dvss.n2510 dvss.n2088 585
R3204 dvss.n2090 dvss.n2089 585
R3205 dvss.n2503 dvss.n2092 585
R3206 dvss.n2502 dvss.n2093 585
R3207 dvss.n2095 dvss.n2094 585
R3208 dvss.n2495 dvss.n2096 585
R3209 dvss.n2494 dvss.n2097 585
R3210 dvss.n2099 dvss.n2098 585
R3211 dvss.n2490 dvss.n2100 585
R3212 dvss.n2489 dvss.n2101 585
R3213 dvss.n2106 dvss.n2102 585
R3214 dvss.n2108 dvss.n2107 585
R3215 dvss.n2482 dvss.n2109 585
R3216 dvss.n2481 dvss.n2110 585
R3217 dvss.n2112 dvss.n2111 585
R3218 dvss.n2477 dvss.n2113 585
R3219 dvss.n2476 dvss.n2114 585
R3220 dvss.n2116 dvss.n2115 585
R3221 dvss.n2472 dvss.n2117 585
R3222 dvss.n2471 dvss.n2118 585
R3223 dvss.n2122 dvss.n2119 585
R3224 dvss.n2464 dvss.n2123 585
R3225 dvss.n2463 dvss.n2124 585
R3226 dvss.n2126 dvss.n2125 585
R3227 dvss.n2456 dvss.n2128 585
R3228 dvss.n2455 dvss.n2129 585
R3229 dvss.n2131 dvss.n2130 585
R3230 dvss.n2448 dvss.n2132 585
R3231 dvss.n2447 dvss.n2133 585
R3232 dvss.n2135 dvss.n2134 585
R3233 dvss.n2443 dvss.n2136 585
R3234 dvss.n2442 dvss.n2137 585
R3235 dvss.n2142 dvss.n2138 585
R3236 dvss.n2144 dvss.n2143 585
R3237 dvss.n2435 dvss.n2145 585
R3238 dvss.n2434 dvss.n2146 585
R3239 dvss.n2148 dvss.n2147 585
R3240 dvss.n2430 dvss.n2149 585
R3241 dvss.n2429 dvss.n2150 585
R3242 dvss.n2152 dvss.n2151 585
R3243 dvss.n2425 dvss.n2153 585
R3244 dvss.n2424 dvss.n2154 585
R3245 dvss.n2158 dvss.n2155 585
R3246 dvss.n2417 dvss.n2159 585
R3247 dvss.n2416 dvss.n2160 585
R3248 dvss.n2162 dvss.n2161 585
R3249 dvss.n2409 dvss.n2164 585
R3250 dvss.n2408 dvss.n2165 585
R3251 dvss.n2167 dvss.n2166 585
R3252 dvss.n2401 dvss.n2168 585
R3253 dvss.n2400 dvss.n2169 585
R3254 dvss.n2171 dvss.n2170 585
R3255 dvss.n2396 dvss.n2172 585
R3256 dvss.n2395 dvss.n2173 585
R3257 dvss.n2178 dvss.n2174 585
R3258 dvss.n2180 dvss.n2179 585
R3259 dvss.n2388 dvss.n2181 585
R3260 dvss.n2387 dvss.n2182 585
R3261 dvss.n2184 dvss.n2183 585
R3262 dvss.n2383 dvss.n2185 585
R3263 dvss.n2382 dvss.n2186 585
R3264 dvss.n2188 dvss.n2187 585
R3265 dvss.n2378 dvss.n2189 585
R3266 dvss.n2377 dvss.n2190 585
R3267 dvss.n2192 dvss.n2191 585
R3268 dvss.n2370 dvss.n1964 585
R3269 dvss.n2666 dvss.n1964 585
R3270 dvss.n2369 dvss.n2195 585
R3271 dvss.n2195 dvss.n1894 585
R3272 dvss.n2218 dvss.n2196 585
R3273 dvss.n2219 dvss.n2218 585
R3274 dvss.n2362 dvss.n2198 585
R3275 dvss.n2220 dvss.n2198 585
R3276 dvss.n2361 dvss.n2199 585
R3277 dvss.n2221 dvss.n2199 585
R3278 dvss.n2222 dvss.n2200 585
R3279 dvss.n2223 dvss.n2222 585
R3280 dvss.n2354 dvss.n2201 585
R3281 dvss.n2225 dvss.n2201 585
R3282 dvss.n2353 dvss.n2202 585
R3283 dvss.n2226 dvss.n2202 585
R3284 dvss.n2227 dvss.n2203 585
R3285 dvss.n2228 dvss.n2227 585
R3286 dvss.n2349 dvss.n2204 585
R3287 dvss.n2229 dvss.n2204 585
R3288 dvss.n2348 dvss.n2205 585
R3289 dvss.n2230 dvss.n2205 585
R3290 dvss.n2232 dvss.n2206 585
R3291 dvss.n2232 dvss.n2231 585
R3292 dvss.n2233 dvss.n2210 585
R3293 dvss.n2234 dvss.n2233 585
R3294 dvss.n2341 dvss.n2211 585
R3295 dvss.n2235 dvss.n2211 585
R3296 dvss.n2340 dvss.n2212 585
R3297 dvss.n2236 dvss.n2212 585
R3298 dvss.n2237 dvss.n2213 585
R3299 dvss.n2238 dvss.n2237 585
R3300 dvss.n2336 dvss.n2214 585
R3301 dvss.n2239 dvss.n2214 585
R3302 dvss.n2335 dvss.n2215 585
R3303 dvss.n2240 dvss.n2215 585
R3304 dvss.n2241 dvss.n2216 585
R3305 dvss.n2242 dvss.n2241 585
R3306 dvss.n2331 dvss.n2217 585
R3307 dvss.n2243 dvss.n2217 585
R3308 dvss.n2330 dvss.n2245 585
R3309 dvss.n2245 dvss.n2244 585
R3310 dvss.n2262 dvss.n2246 585
R3311 dvss.n2263 dvss.n2262 585
R3312 dvss.n2323 dvss.n2249 585
R3313 dvss.n2264 dvss.n2249 585
R3314 dvss.n2322 dvss.n2250 585
R3315 dvss.n2265 dvss.n2250 585
R3316 dvss.n2266 dvss.n2251 585
R3317 dvss.n2267 dvss.n2266 585
R3318 dvss.n2315 dvss.n2253 585
R3319 dvss.n2268 dvss.n2253 585
R3320 dvss.n2314 dvss.n2254 585
R3321 dvss.n2269 dvss.n2254 585
R3322 dvss.n2270 dvss.n2255 585
R3323 dvss.n2271 dvss.n2270 585
R3324 dvss.n2307 dvss.n2256 585
R3325 dvss.n2273 dvss.n2256 585
R3326 dvss.n2306 dvss.n2257 585
R3327 dvss.n2274 dvss.n2257 585
R3328 dvss.n2275 dvss.n2258 585
R3329 dvss.n2276 dvss.n2275 585
R3330 dvss.n2302 dvss.n2259 585
R3331 dvss.n2277 dvss.n2259 585
R3332 dvss.n2301 dvss.n2260 585
R3333 dvss.n2278 dvss.n2260 585
R3334 dvss.n2292 dvss.n2291 585
R3335 dvss.n2291 dvss.n2290 585
R3336 dvss.n2261 dvss.n68 585
R3337 dvss.n2289 dvss.n2261 585
R3338 dvss.n3739 dvss.n69 585
R3339 dvss.n2288 dvss.n69 585
R3340 dvss.n3738 dvss.n70 585
R3341 dvss.n2287 dvss.n70 585
R3342 dvss.n2285 dvss.n71 585
R3343 dvss.n2286 dvss.n2285 585
R3344 dvss.n3734 dvss.n72 585
R3345 dvss.n2284 dvss.n72 585
R3346 dvss.n3733 dvss.n73 585
R3347 dvss.n2283 dvss.n73 585
R3348 dvss.n2281 dvss.n74 585
R3349 dvss.n2282 dvss.n2281 585
R3350 dvss.n3729 dvss.n75 585
R3351 dvss.n2280 dvss.n75 585
R3352 dvss.n3728 dvss.n76 585
R3353 dvss.n2279 dvss.n76 585
R3354 dvss.n1892 dvss.n77 585
R3355 dvss.n1893 dvss.n1892 585
R3356 dvss.n3721 dvss.n80 585
R3357 dvss.n2670 dvss.n80 585
R3358 dvss.n3720 dvss.n81 585
R3359 dvss.n2669 dvss.n81 585
R3360 dvss.n1888 dvss.n82 585
R3361 dvss.n3713 dvss.n84 585
R3362 dvss.n3712 dvss.n85 585
R3363 dvss.n203 dvss.n86 585
R3364 dvss.n204 dvss.n203 585
R3365 dvss.n3705 dvss.n87 585
R3366 dvss.n202 dvss.n87 585
R3367 dvss.n3704 dvss.n88 585
R3368 dvss.n201 dvss.n88 585
R3369 dvss.n199 dvss.n89 585
R3370 dvss.n200 dvss.n199 585
R3371 dvss.n3700 dvss.n90 585
R3372 dvss.n198 dvss.n90 585
R3373 dvss.n3699 dvss.n91 585
R3374 dvss.n197 dvss.n91 585
R3375 dvss.n195 dvss.n92 585
R3376 dvss.n196 dvss.n195 585
R3377 dvss.n194 dvss.n96 585
R3378 dvss.n194 dvss.n193 585
R3379 dvss.n3692 dvss.n97 585
R3380 dvss.n192 dvss.n97 585
R3381 dvss.n3691 dvss.n98 585
R3382 dvss.n191 dvss.n98 585
R3383 dvss.n189 dvss.n99 585
R3384 dvss.n190 dvss.n189 585
R3385 dvss.n3687 dvss.n100 585
R3386 dvss.n188 dvss.n100 585
R3387 dvss.n3686 dvss.n101 585
R3388 dvss.n187 dvss.n101 585
R3389 dvss.n185 dvss.n102 585
R3390 dvss.n186 dvss.n185 585
R3391 dvss.n3682 dvss.n103 585
R3392 dvss.n184 dvss.n103 585
R3393 dvss.n3681 dvss.n104 585
R3394 dvss.n183 dvss.n104 585
R3395 dvss.n181 dvss.n105 585
R3396 dvss.n182 dvss.n181 585
R3397 dvss.n3674 dvss.n108 585
R3398 dvss.n180 dvss.n108 585
R3399 dvss.n3673 dvss.n109 585
R3400 dvss.n179 dvss.n109 585
R3401 dvss.n171 dvss.n110 585
R3402 dvss.n3666 dvss.n112 585
R3403 dvss.n3665 dvss.n113 585
R3404 dvss.n174 dvss.n114 585
R3405 dvss.n175 dvss.n174 585
R3406 dvss.n3658 dvss.n115 585
R3407 dvss.n173 dvss.n115 585
R3408 dvss.n3657 dvss.n116 585
R3409 dvss.n172 dvss.n116 585
R3410 dvss.n118 dvss.n117 585
R3411 dvss.n119 dvss.n118 585
R3412 dvss.n3653 dvss.n3652 585
R3413 dvss.n3652 dvss.n3651 585
R3414 dvss.n3650 dvss.n3649 583.256
R3415 dvss.n3442 dvss.n3439 564.282
R3416 dvss.n3264 dvss.n259 564.282
R3417 dvss.n3148 dvss.n323 564.282
R3418 dvss.n3023 dvss.n3021 564.282
R3419 dvss.n2895 dvss.n447 564.282
R3420 dvss.n1480 dvss.n1477 564.282
R3421 dvss.n1306 dvss.n556 564.282
R3422 dvss.n717 dvss.n626 564.282
R3423 dvss.n899 dvss.n877 539.294
R3424 dvss.n895 dvss.n877 539.294
R3425 dvss.n895 dvss.n881 539.294
R3426 dvss.n891 dvss.n881 539.294
R3427 dvss.n891 dvss.n883 539.294
R3428 dvss.n883 dvss.n874 539.294
R3429 dvss.n907 dvss.n874 539.294
R3430 dvss.n907 dvss.n871 539.294
R3431 dvss.n921 dvss.n871 539.294
R3432 dvss.n921 dvss.n870 539.294
R3433 dvss.n926 dvss.n870 539.294
R3434 dvss.n926 dvss.n866 539.294
R3435 dvss.n940 dvss.n866 539.294
R3436 dvss.n940 dvss.n864 539.294
R3437 dvss.n944 dvss.n864 539.294
R3438 dvss.n945 dvss.n944 539.294
R3439 dvss.n947 dvss.n764 539.294
R3440 dvss.n960 dvss.n764 539.294
R3441 dvss.n960 dvss.n759 539.294
R3442 dvss.n969 dvss.n759 539.294
R3443 dvss.n970 dvss.n969 539.294
R3444 dvss.n970 dvss.n749 539.294
R3445 dvss.n983 dvss.n749 539.294
R3446 dvss.n989 dvss.n983 539.294
R3447 dvss.n989 dvss.n988 539.294
R3448 dvss.n988 dvss.n739 539.294
R3449 dvss.n1006 dvss.n739 539.294
R3450 dvss.n1006 dvss.n731 539.294
R3451 dvss.n1021 dvss.n731 539.294
R3452 dvss.n1022 dvss.n1021 539.294
R3453 dvss.n1022 dvss.n730 539.294
R3454 dvss.n1027 dvss.n730 539.294
R3455 dvss.n1027 dvss.n617 539.294
R3456 dvss.n1106 dvss.n617 539.294
R3457 dvss.n1106 dvss.n618 539.294
R3458 dvss.n1102 dvss.n618 539.294
R3459 dvss.n1050 dvss.n624 539.294
R3460 dvss.n1097 dvss.n628 539.294
R3461 dvss.n1097 dvss.n629 539.294
R3462 dvss.n1093 dvss.n629 539.294
R3463 dvss.n1093 dvss.n635 539.294
R3464 dvss.n1089 dvss.n635 539.294
R3465 dvss.n1089 dvss.n639 539.294
R3466 dvss.n1085 dvss.n639 539.294
R3467 dvss.n1085 dvss.n644 539.294
R3468 dvss.n671 dvss.n644 539.294
R3469 dvss.n678 dvss.n671 539.294
R3470 dvss.n679 dvss.n678 539.294
R3471 dvss.n679 dvss.n668 539.294
R3472 dvss.n685 dvss.n668 539.294
R3473 dvss.n686 dvss.n685 539.294
R3474 dvss.n686 dvss.n569 539.294
R3475 dvss.n1294 dvss.n569 539.294
R3476 dvss.n1294 dvss.n560 539.294
R3477 dvss.n1321 dvss.n560 539.294
R3478 dvss.n1321 dvss.n561 539.294
R3479 dvss.n1310 dvss.n561 539.294
R3480 dvss.n1312 dvss.n1309 539.294
R3481 dvss.n1309 dvss.n550 539.294
R3482 dvss.n1336 dvss.n550 539.294
R3483 dvss.n1336 dvss.n546 539.294
R3484 dvss.n1349 dvss.n546 539.294
R3485 dvss.n1350 dvss.n1349 539.294
R3486 dvss.n1350 dvss.n540 539.294
R3487 dvss.n540 dvss.n535 539.294
R3488 dvss.n1373 dvss.n535 539.294
R3489 dvss.n1374 dvss.n1373 539.294
R3490 dvss.n1374 dvss.n531 539.294
R3491 dvss.n531 dvss.n525 539.294
R3492 dvss.n1398 dvss.n525 539.294
R3493 dvss.n1399 dvss.n1398 539.294
R3494 dvss.n1399 dvss.n524 539.294
R3495 dvss.n1404 dvss.n524 539.294
R3496 dvss.n1404 dvss.n507 539.294
R3497 dvss.n1579 dvss.n507 539.294
R3498 dvss.n1579 dvss.n508 539.294
R3499 dvss.n1486 dvss.n508 539.294
R3500 dvss.n1485 dvss.n1484 539.294
R3501 dvss.n1492 dvss.n1490 539.294
R3502 dvss.n1492 dvss.n1475 539.294
R3503 dvss.n1496 dvss.n1475 539.294
R3504 dvss.n1497 dvss.n1496 539.294
R3505 dvss.n1502 dvss.n1497 539.294
R3506 dvss.n1502 dvss.n1471 539.294
R3507 dvss.n1507 dvss.n1471 539.294
R3508 dvss.n1508 dvss.n1507 539.294
R3509 dvss.n1508 dvss.n1469 539.294
R3510 dvss.n1515 dvss.n1469 539.294
R3511 dvss.n1516 dvss.n1515 539.294
R3512 dvss.n1516 dvss.n1466 539.294
R3513 dvss.n1522 dvss.n1466 539.294
R3514 dvss.n1523 dvss.n1522 539.294
R3515 dvss.n1523 dvss.n459 539.294
R3516 dvss.n2884 dvss.n459 539.294
R3517 dvss.n2884 dvss.n451 539.294
R3518 dvss.n2913 dvss.n451 539.294
R3519 dvss.n2913 dvss.n452 539.294
R3520 dvss.n2904 dvss.n2901 539.294
R3521 dvss.n2902 dvss.n441 539.294
R3522 dvss.n2928 dvss.n441 539.294
R3523 dvss.n2928 dvss.n437 539.294
R3524 dvss.n2941 dvss.n437 539.294
R3525 dvss.n2942 dvss.n2941 539.294
R3526 dvss.n2942 dvss.n431 539.294
R3527 dvss.n431 dvss.n426 539.294
R3528 dvss.n2965 dvss.n426 539.294
R3529 dvss.n2966 dvss.n2965 539.294
R3530 dvss.n2966 dvss.n422 539.294
R3531 dvss.n422 dvss.n416 539.294
R3532 dvss.n2990 dvss.n416 539.294
R3533 dvss.n2991 dvss.n2990 539.294
R3534 dvss.n2991 dvss.n415 539.294
R3535 dvss.n2997 dvss.n415 539.294
R3536 dvss.n2997 dvss.n399 539.294
R3537 dvss.n3014 dvss.n399 539.294
R3538 dvss.n3014 dvss.n393 539.294
R3539 dvss.n3033 dvss.n393 539.294
R3540 dvss.n392 dvss.n389 539.294
R3541 dvss.n3037 dvss.n382 539.294
R3542 dvss.n3050 dvss.n382 539.294
R3543 dvss.n3050 dvss.n379 539.294
R3544 dvss.n3057 dvss.n379 539.294
R3545 dvss.n3057 dvss.n372 539.294
R3546 dvss.n3076 dvss.n372 539.294
R3547 dvss.n3076 dvss.n367 539.294
R3548 dvss.n3081 dvss.n367 539.294
R3549 dvss.n3081 dvss.n361 539.294
R3550 dvss.n3093 dvss.n361 539.294
R3551 dvss.n3093 dvss.n356 539.294
R3552 dvss.n3107 dvss.n356 539.294
R3553 dvss.n3107 dvss.n352 539.294
R3554 dvss.n3114 dvss.n352 539.294
R3555 dvss.n3114 dvss.n353 539.294
R3556 dvss.n353 dvss.n341 539.294
R3557 dvss.n341 dvss.n334 539.294
R3558 dvss.n3135 dvss.n334 539.294
R3559 dvss.n3136 dvss.n3135 539.294
R3560 dvss.n3140 dvss.n330 539.294
R3561 dvss.n331 dvss.n317 539.294
R3562 dvss.n3167 dvss.n317 539.294
R3563 dvss.n3167 dvss.n314 539.294
R3564 dvss.n3174 dvss.n314 539.294
R3565 dvss.n3174 dvss.n307 539.294
R3566 dvss.n3189 dvss.n307 539.294
R3567 dvss.n3189 dvss.n303 539.294
R3568 dvss.n3197 dvss.n303 539.294
R3569 dvss.n3197 dvss.n297 539.294
R3570 dvss.n3209 dvss.n297 539.294
R3571 dvss.n3209 dvss.n292 539.294
R3572 dvss.n3223 dvss.n292 539.294
R3573 dvss.n3223 dvss.n288 539.294
R3574 dvss.n3230 dvss.n288 539.294
R3575 dvss.n3230 dvss.n289 539.294
R3576 dvss.n289 dvss.n277 539.294
R3577 dvss.n277 dvss.n270 539.294
R3578 dvss.n3251 dvss.n270 539.294
R3579 dvss.n3252 dvss.n3251 539.294
R3580 dvss.n3256 dvss.n266 539.294
R3581 dvss.n267 dvss.n256 539.294
R3582 dvss.n256 dvss.n251 539.294
R3583 dvss.n3288 dvss.n251 539.294
R3584 dvss.n3289 dvss.n3288 539.294
R3585 dvss.n3289 dvss.n240 539.294
R3586 dvss.n3308 dvss.n240 539.294
R3587 dvss.n3308 dvss.n236 539.294
R3588 dvss.n3313 dvss.n236 539.294
R3589 dvss.n3314 dvss.n3313 539.294
R3590 dvss.n3314 dvss.n232 539.294
R3591 dvss.n232 dvss.n226 539.294
R3592 dvss.n3338 dvss.n226 539.294
R3593 dvss.n3339 dvss.n3338 539.294
R3594 dvss.n3339 dvss.n225 539.294
R3595 dvss.n3344 dvss.n225 539.294
R3596 dvss.n3344 dvss.n208 539.294
R3597 dvss.n3545 dvss.n208 539.294
R3598 dvss.n3545 dvss.n209 539.294
R3599 dvss.n3435 dvss.n209 539.294
R3600 dvss.n3434 dvss.n3433 539.294
R3601 dvss.n3431 dvss.n3430 539.294
R3602 dvss.n3448 dvss.n3430 539.294
R3603 dvss.n3449 dvss.n3448 539.294
R3604 dvss.n3449 dvss.n3424 539.294
R3605 dvss.n3455 dvss.n3424 539.294
R3606 dvss.n3457 dvss.n3455 539.294
R3607 dvss.n3457 dvss.n3456 539.294
R3608 dvss.n3456 dvss.n3421 539.294
R3609 dvss.n3465 dvss.n3421 539.294
R3610 dvss.n3467 dvss.n3465 539.294
R3611 dvss.n3468 dvss.n3467 539.294
R3612 dvss.n3469 dvss.n3468 539.294
R3613 dvss.n3469 dvss.n3414 539.294
R3614 dvss.n3477 dvss.n3414 539.294
R3615 dvss.n3477 dvss.n3410 539.294
R3616 dvss.n3483 dvss.n3410 539.294
R3617 dvss.n3484 dvss.n3483 539.294
R3618 dvss.n3487 dvss.n3484 539.294
R3619 dvss.n3488 dvss.n3487 539.294
R3620 dvss.n3488 dvss.n122 539.294
R3621 dvss.n851 dvss.n766 539.294
R3622 dvss.n851 dvss.n850 539.294
R3623 dvss.n850 dvss.n772 539.294
R3624 dvss.n846 dvss.n772 539.294
R3625 dvss.n846 dvss.n774 539.294
R3626 dvss.n842 dvss.n774 539.294
R3627 dvss.n842 dvss.n780 539.294
R3628 dvss.n838 dvss.n780 539.294
R3629 dvss.n838 dvss.n781 539.294
R3630 dvss.n834 dvss.n781 539.294
R3631 dvss.n834 dvss.n805 539.294
R3632 dvss.n830 dvss.n805 539.294
R3633 dvss.n830 dvss.n807 539.294
R3634 dvss.n826 dvss.n807 539.294
R3635 dvss.n826 dvss.n822 539.294
R3636 dvss.n822 dvss.n612 539.294
R3637 dvss.n1112 dvss.n612 539.294
R3638 dvss.n1112 dvss.n609 539.294
R3639 dvss.n1119 dvss.n609 539.294
R3640 dvss.n1123 dvss.n608 539.294
R3641 dvss.n1131 dvss.n605 539.294
R3642 dvss.n1131 dvss.n603 539.294
R3643 dvss.n1135 dvss.n603 539.294
R3644 dvss.n1135 dvss.n597 539.294
R3645 dvss.n1146 dvss.n597 539.294
R3646 dvss.n1146 dvss.n595 539.294
R3647 dvss.n1151 dvss.n595 539.294
R3648 dvss.n1151 dvss.n587 539.294
R3649 dvss.n1161 dvss.n587 539.294
R3650 dvss.n1161 dvss.n586 539.294
R3651 dvss.n1166 dvss.n586 539.294
R3652 dvss.n1166 dvss.n579 539.294
R3653 dvss.n1176 dvss.n579 539.294
R3654 dvss.n1176 dvss.n578 539.294
R3655 dvss.n1180 dvss.n578 539.294
R3656 dvss.n1180 dvss.n573 539.294
R3657 dvss.n1289 dvss.n573 539.294
R3658 dvss.n1289 dvss.n574 539.294
R3659 dvss.n1184 dvss.n574 539.294
R3660 dvss.n1212 dvss.n1185 539.294
R3661 dvss.n1188 dvss.n1187 539.294
R3662 dvss.n1219 dvss.n1188 539.294
R3663 dvss.n1220 dvss.n1219 539.294
R3664 dvss.n1220 dvss.n1193 539.294
R3665 dvss.n1194 dvss.n1193 539.294
R3666 dvss.n1211 dvss.n1194 539.294
R3667 dvss.n1211 dvss.n1199 539.294
R3668 dvss.n1200 dvss.n1199 539.294
R3669 dvss.n1229 dvss.n1200 539.294
R3670 dvss.n1229 dvss.n1203 539.294
R3671 dvss.n1204 dvss.n1203 539.294
R3672 dvss.n1234 dvss.n1204 539.294
R3673 dvss.n1235 dvss.n1234 539.294
R3674 dvss.n1235 dvss.n1210 539.294
R3675 dvss.n1239 dvss.n1210 539.294
R3676 dvss.n1239 dvss.n502 539.294
R3677 dvss.n1585 dvss.n502 539.294
R3678 dvss.n1585 dvss.n499 539.294
R3679 dvss.n1592 dvss.n499 539.294
R3680 dvss.n1596 dvss.n498 539.294
R3681 dvss.n1604 dvss.n495 539.294
R3682 dvss.n1604 dvss.n493 539.294
R3683 dvss.n1608 dvss.n493 539.294
R3684 dvss.n1608 dvss.n487 539.294
R3685 dvss.n1619 dvss.n487 539.294
R3686 dvss.n1619 dvss.n485 539.294
R3687 dvss.n1624 dvss.n485 539.294
R3688 dvss.n1624 dvss.n477 539.294
R3689 dvss.n1634 dvss.n477 539.294
R3690 dvss.n1634 dvss.n476 539.294
R3691 dvss.n1639 dvss.n476 539.294
R3692 dvss.n1639 dvss.n469 539.294
R3693 dvss.n1649 dvss.n469 539.294
R3694 dvss.n1649 dvss.n468 539.294
R3695 dvss.n1653 dvss.n468 539.294
R3696 dvss.n1653 dvss.n463 539.294
R3697 dvss.n2879 dvss.n463 539.294
R3698 dvss.n2879 dvss.n464 539.294
R3699 dvss.n1657 dvss.n464 539.294
R3700 dvss.n1792 dvss.n1658 539.294
R3701 dvss.n1661 dvss.n1660 539.294
R3702 dvss.n1799 dvss.n1661 539.294
R3703 dvss.n1800 dvss.n1799 539.294
R3704 dvss.n1800 dvss.n1666 539.294
R3705 dvss.n1667 dvss.n1666 539.294
R3706 dvss.n1791 dvss.n1667 539.294
R3707 dvss.n1791 dvss.n1672 539.294
R3708 dvss.n1673 dvss.n1672 539.294
R3709 dvss.n1809 dvss.n1673 539.294
R3710 dvss.n1809 dvss.n1676 539.294
R3711 dvss.n1677 dvss.n1676 539.294
R3712 dvss.n1814 dvss.n1677 539.294
R3713 dvss.n1815 dvss.n1814 539.294
R3714 dvss.n1815 dvss.n1683 539.294
R3715 dvss.n1684 dvss.n1683 539.294
R3716 dvss.n1819 dvss.n1684 539.294
R3717 dvss.n1819 dvss.n1686 539.294
R3718 dvss.n1687 dvss.n1686 539.294
R3719 dvss.n1788 dvss.n1687 539.294
R3720 dvss.n1690 dvss.n1689 539.294
R3721 dvss.n1786 dvss.n1692 539.294
R3722 dvss.n1693 dvss.n1692 539.294
R3723 dvss.n1827 dvss.n1693 539.294
R3724 dvss.n1827 dvss.n1697 539.294
R3725 dvss.n1698 dvss.n1697 539.294
R3726 dvss.n1785 dvss.n1698 539.294
R3727 dvss.n1785 dvss.n1703 539.294
R3728 dvss.n1704 dvss.n1703 539.294
R3729 dvss.n1834 dvss.n1704 539.294
R3730 dvss.n1834 dvss.n1707 539.294
R3731 dvss.n1708 dvss.n1707 539.294
R3732 dvss.n1839 dvss.n1708 539.294
R3733 dvss.n1840 dvss.n1839 539.294
R3734 dvss.n1840 dvss.n1714 539.294
R3735 dvss.n1715 dvss.n1714 539.294
R3736 dvss.n1844 dvss.n1715 539.294
R3737 dvss.n1844 dvss.n1717 539.294
R3738 dvss.n1718 dvss.n1717 539.294
R3739 dvss.n1782 dvss.n1718 539.294
R3740 dvss.n1721 dvss.n1720 539.294
R3741 dvss.n1780 dvss.n1723 539.294
R3742 dvss.n1724 dvss.n1723 539.294
R3743 dvss.n1852 dvss.n1724 539.294
R3744 dvss.n1852 dvss.n1728 539.294
R3745 dvss.n1729 dvss.n1728 539.294
R3746 dvss.n1779 dvss.n1729 539.294
R3747 dvss.n1779 dvss.n1734 539.294
R3748 dvss.n1735 dvss.n1734 539.294
R3749 dvss.n1859 dvss.n1735 539.294
R3750 dvss.n1859 dvss.n1738 539.294
R3751 dvss.n1739 dvss.n1738 539.294
R3752 dvss.n1864 dvss.n1739 539.294
R3753 dvss.n1865 dvss.n1864 539.294
R3754 dvss.n1865 dvss.n1745 539.294
R3755 dvss.n1746 dvss.n1745 539.294
R3756 dvss.n1869 dvss.n1746 539.294
R3757 dvss.n1869 dvss.n1748 539.294
R3758 dvss.n1749 dvss.n1748 539.294
R3759 dvss.n1876 dvss.n1749 539.294
R3760 dvss.n1752 dvss.n1751 539.294
R3761 dvss.n1874 dvss.n1754 539.294
R3762 dvss.n1755 dvss.n1754 539.294
R3763 dvss.n1882 dvss.n1755 539.294
R3764 dvss.n1882 dvss.n1759 539.294
R3765 dvss.n1760 dvss.n1759 539.294
R3766 dvss.n1778 dvss.n1760 539.294
R3767 dvss.n1778 dvss.n1765 539.294
R3768 dvss.n1766 dvss.n1765 539.294
R3769 dvss.n2674 dvss.n1766 539.294
R3770 dvss.n2674 dvss.n1769 539.294
R3771 dvss.n1770 dvss.n1769 539.294
R3772 dvss.n2678 dvss.n1770 539.294
R3773 dvss.n2678 dvss.n1777 539.294
R3774 dvss.n2682 dvss.n1777 539.294
R3775 dvss.n2682 dvss.n169 539.294
R3776 dvss.n3550 dvss.n169 539.294
R3777 dvss.n3550 dvss.n164 539.294
R3778 dvss.n3569 dvss.n164 539.294
R3779 dvss.n3569 dvss.n165 539.294
R3780 dvss.n3556 dvss.n3555 539.294
R3781 dvss.n3558 dvss.n161 539.294
R3782 dvss.n3575 dvss.n161 539.294
R3783 dvss.n3575 dvss.n156 539.294
R3784 dvss.n3588 dvss.n156 539.294
R3785 dvss.n3588 dvss.n155 539.294
R3786 dvss.n3592 dvss.n155 539.294
R3787 dvss.n3592 dvss.n148 539.294
R3788 dvss.n3603 dvss.n148 539.294
R3789 dvss.n3603 dvss.n145 539.294
R3790 dvss.n3607 dvss.n145 539.294
R3791 dvss.n3607 dvss.n142 539.294
R3792 dvss.n3621 dvss.n142 539.294
R3793 dvss.n3621 dvss.n140 539.294
R3794 dvss.n3625 dvss.n140 539.294
R3795 dvss.n3625 dvss.n136 539.294
R3796 dvss.n3634 dvss.n136 539.294
R3797 dvss.n3634 dvss.n132 539.294
R3798 dvss.n3639 dvss.n132 539.294
R3799 dvss.n3640 dvss.n3639 539.294
R3800 dvss.n958 dvss.n858 539.294
R3801 dvss.n958 dvss.n760 539.294
R3802 dvss.n967 dvss.n760 539.294
R3803 dvss.n967 dvss.n752 539.294
R3804 dvss.n980 dvss.n752 539.294
R3805 dvss.n980 dvss.n747 539.294
R3806 dvss.n991 dvss.n747 539.294
R3807 dvss.n991 dvss.n740 539.294
R3808 dvss.n1002 dvss.n740 539.294
R3809 dvss.n1002 dvss.n734 539.294
R3810 dvss.n1018 dvss.n734 539.294
R3811 dvss.n1019 dvss.n1018 539.294
R3812 dvss.n1019 dvss.n727 539.294
R3813 dvss.n728 dvss.n727 539.294
R3814 dvss.n1025 dvss.n728 539.294
R3815 dvss.n1025 dvss.n719 539.294
R3816 dvss.n719 dvss.n615 539.294
R3817 dvss.n1044 dvss.n615 539.294
R3818 dvss.n1045 dvss.n1044 539.294
R3819 dvss.n1047 dvss.n715 539.294
R3820 dvss.n713 dvss.n627 539.294
R3821 dvss.n1062 dvss.n627 539.294
R3822 dvss.n1062 dvss.n636 539.294
R3823 dvss.n637 dvss.n636 539.294
R3824 dvss.n638 dvss.n637 539.294
R3825 dvss.n647 dvss.n638 539.294
R3826 dvss.n1083 dvss.n647 539.294
R3827 dvss.n1083 dvss.n648 539.294
R3828 dvss.n674 dvss.n648 539.294
R3829 dvss.n674 dvss.n654 539.294
R3830 dvss.n655 dvss.n654 539.294
R3831 dvss.n682 dvss.n655 539.294
R3832 dvss.n683 dvss.n682 539.294
R3833 dvss.n683 dvss.n667 539.294
R3834 dvss.n689 dvss.n667 539.294
R3835 dvss.n689 dvss.n570 539.294
R3836 dvss.n570 dvss.n566 539.294
R3837 dvss.n566 dvss.n559 539.294
R3838 dvss.n1303 dvss.n559 539.294
R3839 dvss.n1308 dvss.n1304 539.294
R3840 dvss.n1325 dvss.n555 539.294
R3841 dvss.n1325 dvss.n549 539.294
R3842 dvss.n1339 dvss.n549 539.294
R3843 dvss.n1339 dvss.n543 539.294
R3844 dvss.n1352 dvss.n543 539.294
R3845 dvss.n1352 dvss.n537 539.294
R3846 dvss.n1368 dvss.n537 539.294
R3847 dvss.n1368 dvss.n534 539.294
R3848 dvss.n1376 dvss.n534 539.294
R3849 dvss.n1376 dvss.n528 539.294
R3850 dvss.n1395 dvss.n528 539.294
R3851 dvss.n1396 dvss.n1395 539.294
R3852 dvss.n1396 dvss.n521 539.294
R3853 dvss.n522 dvss.n521 539.294
R3854 dvss.n1402 dvss.n522 539.294
R3855 dvss.n1402 dvss.n513 539.294
R3856 dvss.n513 dvss.n505 539.294
R3857 dvss.n1418 dvss.n505 539.294
R3858 dvss.n1478 dvss.n1418 539.294
R3859 dvss.n1423 dvss.n1422 539.294
R3860 dvss.n1483 dvss.n1482 539.294
R3861 dvss.n1483 dvss.n1432 539.294
R3862 dvss.n1433 dvss.n1432 539.294
R3863 dvss.n1473 dvss.n1433 539.294
R3864 dvss.n1474 dvss.n1473 539.294
R3865 dvss.n1474 dvss.n1443 539.294
R3866 dvss.n1444 dvss.n1443 539.294
R3867 dvss.n1510 dvss.n1444 539.294
R3868 dvss.n1511 dvss.n1510 539.294
R3869 dvss.n1511 dvss.n1452 539.294
R3870 dvss.n1453 dvss.n1452 539.294
R3871 dvss.n1519 dvss.n1453 539.294
R3872 dvss.n1520 dvss.n1519 539.294
R3873 dvss.n1520 dvss.n1465 539.294
R3874 dvss.n1526 dvss.n1465 539.294
R3875 dvss.n1526 dvss.n460 539.294
R3876 dvss.n460 dvss.n456 539.294
R3877 dvss.n456 dvss.n450 539.294
R3878 dvss.n2892 dvss.n450 539.294
R3879 dvss.n2897 dvss.n2893 539.294
R3880 dvss.n2917 dvss.n446 539.294
R3881 dvss.n2917 dvss.n440 539.294
R3882 dvss.n2931 dvss.n440 539.294
R3883 dvss.n2931 dvss.n434 539.294
R3884 dvss.n2944 dvss.n434 539.294
R3885 dvss.n2944 dvss.n428 539.294
R3886 dvss.n2960 dvss.n428 539.294
R3887 dvss.n2960 dvss.n425 539.294
R3888 dvss.n2968 dvss.n425 539.294
R3889 dvss.n2968 dvss.n419 539.294
R3890 dvss.n2987 dvss.n419 539.294
R3891 dvss.n2988 dvss.n2987 539.294
R3892 dvss.n2988 dvss.n412 539.294
R3893 dvss.n413 dvss.n412 539.294
R3894 dvss.n2994 dvss.n413 539.294
R3895 dvss.n2994 dvss.n404 539.294
R3896 dvss.n404 dvss.n397 539.294
R3897 dvss.n3017 dvss.n397 539.294
R3898 dvss.n3018 dvss.n3017 539.294
R3899 dvss.n3025 dvss.n3019 539.294
R3900 dvss.n3020 dvss.n387 539.294
R3901 dvss.n387 dvss.n380 539.294
R3902 dvss.n3053 dvss.n380 539.294
R3903 dvss.n3054 dvss.n3053 539.294
R3904 dvss.n3054 dvss.n375 539.294
R3905 dvss.n375 dvss.n371 539.294
R3906 dvss.n371 dvss.n370 539.294
R3907 dvss.n370 dvss.n365 539.294
R3908 dvss.n365 dvss.n359 539.294
R3909 dvss.n3095 dvss.n359 539.294
R3910 dvss.n3096 dvss.n3095 539.294
R3911 dvss.n3096 dvss.n355 539.294
R3912 dvss.n355 dvss.n349 539.294
R3913 dvss.n350 dvss.n349 539.294
R3914 dvss.n3110 dvss.n350 539.294
R3915 dvss.n3110 dvss.n337 539.294
R3916 dvss.n3132 dvss.n337 539.294
R3917 dvss.n3132 dvss.n325 539.294
R3918 dvss.n3146 dvss.n325 539.294
R3919 dvss.n324 dvss.n322 539.294
R3920 dvss.n3150 dvss.n315 539.294
R3921 dvss.n3169 dvss.n315 539.294
R3922 dvss.n3170 dvss.n3169 539.294
R3923 dvss.n3170 dvss.n312 539.294
R3924 dvss.n312 dvss.n305 539.294
R3925 dvss.n3191 dvss.n305 539.294
R3926 dvss.n3192 dvss.n3191 539.294
R3927 dvss.n3192 dvss.n301 539.294
R3928 dvss.n301 dvss.n295 539.294
R3929 dvss.n3211 dvss.n295 539.294
R3930 dvss.n3212 dvss.n3211 539.294
R3931 dvss.n3212 dvss.n291 539.294
R3932 dvss.n291 dvss.n285 539.294
R3933 dvss.n286 dvss.n285 539.294
R3934 dvss.n3226 dvss.n286 539.294
R3935 dvss.n3226 dvss.n273 539.294
R3936 dvss.n3248 dvss.n273 539.294
R3937 dvss.n3248 dvss.n261 539.294
R3938 dvss.n3262 dvss.n261 539.294
R3939 dvss.n260 dvss.n258 539.294
R3940 dvss.n3266 dvss.n253 539.294
R3941 dvss.n3285 dvss.n253 539.294
R3942 dvss.n3285 dvss.n248 539.294
R3943 dvss.n3291 dvss.n248 539.294
R3944 dvss.n3291 dvss.n249 539.294
R3945 dvss.n249 dvss.n239 539.294
R3946 dvss.n244 dvss.n239 539.294
R3947 dvss.n244 dvss.n235 539.294
R3948 dvss.n3316 dvss.n235 539.294
R3949 dvss.n3316 dvss.n229 539.294
R3950 dvss.n3335 dvss.n229 539.294
R3951 dvss.n3336 dvss.n3335 539.294
R3952 dvss.n3336 dvss.n222 539.294
R3953 dvss.n223 dvss.n222 539.294
R3954 dvss.n3342 dvss.n223 539.294
R3955 dvss.n3342 dvss.n214 539.294
R3956 dvss.n214 dvss.n206 539.294
R3957 dvss.n3358 dvss.n206 539.294
R3958 dvss.n3440 dvss.n3358 539.294
R3959 dvss.n3363 dvss.n3362 539.294
R3960 dvss.n3445 dvss.n3444 539.294
R3961 dvss.n3445 dvss.n3372 539.294
R3962 dvss.n3373 dvss.n3372 539.294
R3963 dvss.n3452 dvss.n3373 539.294
R3964 dvss.n3453 dvss.n3452 539.294
R3965 dvss.n3453 dvss.n3383 539.294
R3966 dvss.n3384 dvss.n3383 539.294
R3967 dvss.n3462 dvss.n3384 539.294
R3968 dvss.n3463 dvss.n3462 539.294
R3969 dvss.n3463 dvss.n3392 539.294
R3970 dvss.n3393 dvss.n3392 539.294
R3971 dvss.n3419 dvss.n3393 539.294
R3972 dvss.n3472 dvss.n3419 539.294
R3973 dvss.n3472 dvss.n3412 539.294
R3974 dvss.n3480 dvss.n3412 539.294
R3975 dvss.n3481 dvss.n3480 539.294
R3976 dvss.n3481 dvss.n3407 539.294
R3977 dvss.n3408 dvss.n3407 539.294
R3978 dvss.n3408 dvss.n123 539.294
R3979 dvss.n3648 dvss.n123 539.294
R3980 dvss.n2665 dvss.n1965 539.294
R3981 dvss.n1968 dvss.n1967 539.294
R3982 dvss.n1971 dvss.n1970 539.294
R3983 dvss.n1973 dvss.n1972 539.294
R3984 dvss.n1976 dvss.n1975 539.294
R3985 dvss.n1982 dvss.n1981 539.294
R3986 dvss.n1984 dvss.n1983 539.294
R3987 dvss.n1992 dvss.n1991 539.294
R3988 dvss.n1994 dvss.n1993 539.294
R3989 dvss.n1996 dvss.n1995 539.294
R3990 dvss.n2002 dvss.n2001 539.294
R3991 dvss.n2005 dvss.n2004 539.294
R3992 dvss.n2007 dvss.n2006 539.294
R3993 dvss.n2010 dvss.n2009 539.294
R3994 dvss.n2015 dvss.n2014 539.294
R3995 dvss.n2017 dvss.n2016 539.294
R3996 dvss.n2021 dvss.n2020 539.294
R3997 dvss.n2024 dvss.n2023 539.294
R3998 dvss.n2026 dvss.n2025 539.294
R3999 dvss.n2029 dvss.n2028 539.294
R4000 dvss.n2035 dvss.n2034 539.294
R4001 dvss.n2038 dvss.n2037 539.294
R4002 dvss.n2041 dvss.n2040 539.294
R4003 dvss.n2043 dvss.n2042 539.294
R4004 dvss.n2046 dvss.n2045 539.294
R4005 dvss.n2051 dvss.n2050 539.294
R4006 dvss.n2053 dvss.n2052 539.294
R4007 dvss.n2057 dvss.n2056 539.294
R4008 dvss.n2060 dvss.n2059 539.294
R4009 dvss.n2062 dvss.n2061 539.294
R4010 dvss.n2065 dvss.n2064 539.294
R4011 dvss.n2071 dvss.n2070 539.294
R4012 dvss.n2074 dvss.n2073 539.294
R4013 dvss.n2077 dvss.n2076 539.294
R4014 dvss.n2079 dvss.n2078 539.294
R4015 dvss.n2082 dvss.n2081 539.294
R4016 dvss.n2087 dvss.n2086 539.294
R4017 dvss.n2089 dvss.n2088 539.294
R4018 dvss.n2093 dvss.n2092 539.294
R4019 dvss.n2096 dvss.n2095 539.294
R4020 dvss.n2098 dvss.n2097 539.294
R4021 dvss.n2101 dvss.n2100 539.294
R4022 dvss.n2107 dvss.n2106 539.294
R4023 dvss.n2110 dvss.n2109 539.294
R4024 dvss.n2113 dvss.n2112 539.294
R4025 dvss.n2115 dvss.n2114 539.294
R4026 dvss.n2118 dvss.n2117 539.294
R4027 dvss.n2123 dvss.n2122 539.294
R4028 dvss.n2125 dvss.n2124 539.294
R4029 dvss.n2129 dvss.n2128 539.294
R4030 dvss.n2132 dvss.n2131 539.294
R4031 dvss.n2134 dvss.n2133 539.294
R4032 dvss.n2137 dvss.n2136 539.294
R4033 dvss.n2143 dvss.n2142 539.294
R4034 dvss.n2146 dvss.n2145 539.294
R4035 dvss.n2149 dvss.n2148 539.294
R4036 dvss.n2151 dvss.n2150 539.294
R4037 dvss.n2154 dvss.n2153 539.294
R4038 dvss.n2159 dvss.n2158 539.294
R4039 dvss.n2161 dvss.n2160 539.294
R4040 dvss.n2165 dvss.n2164 539.294
R4041 dvss.n2168 dvss.n2167 539.294
R4042 dvss.n2170 dvss.n2169 539.294
R4043 dvss.n2173 dvss.n2172 539.294
R4044 dvss.n2179 dvss.n2178 539.294
R4045 dvss.n2182 dvss.n2181 539.294
R4046 dvss.n2185 dvss.n2184 539.294
R4047 dvss.n2187 dvss.n2186 539.294
R4048 dvss.n2190 dvss.n2189 539.294
R4049 dvss.n2191 dvss.n1964 539.294
R4050 dvss.n2195 dvss.n1964 539.294
R4051 dvss.n2218 dvss.n2195 539.294
R4052 dvss.n2218 dvss.n2198 539.294
R4053 dvss.n2199 dvss.n2198 539.294
R4054 dvss.n2222 dvss.n2199 539.294
R4055 dvss.n2222 dvss.n2201 539.294
R4056 dvss.n2202 dvss.n2201 539.294
R4057 dvss.n2227 dvss.n2202 539.294
R4058 dvss.n2227 dvss.n2204 539.294
R4059 dvss.n2205 dvss.n2204 539.294
R4060 dvss.n2232 dvss.n2205 539.294
R4061 dvss.n2233 dvss.n2232 539.294
R4062 dvss.n2233 dvss.n2211 539.294
R4063 dvss.n2212 dvss.n2211 539.294
R4064 dvss.n2237 dvss.n2212 539.294
R4065 dvss.n2237 dvss.n2214 539.294
R4066 dvss.n2215 dvss.n2214 539.294
R4067 dvss.n2241 dvss.n2215 539.294
R4068 dvss.n2241 dvss.n2217 539.294
R4069 dvss.n2245 dvss.n2217 539.294
R4070 dvss.n2262 dvss.n2245 539.294
R4071 dvss.n2262 dvss.n2249 539.294
R4072 dvss.n2250 dvss.n2249 539.294
R4073 dvss.n2266 dvss.n2250 539.294
R4074 dvss.n2266 dvss.n2253 539.294
R4075 dvss.n2254 dvss.n2253 539.294
R4076 dvss.n2270 dvss.n2254 539.294
R4077 dvss.n2270 dvss.n2256 539.294
R4078 dvss.n2257 dvss.n2256 539.294
R4079 dvss.n2275 dvss.n2257 539.294
R4080 dvss.n2275 dvss.n2259 539.294
R4081 dvss.n2260 dvss.n2259 539.294
R4082 dvss.n2291 dvss.n2260 539.294
R4083 dvss.n2291 dvss.n2261 539.294
R4084 dvss.n2261 dvss.n69 539.294
R4085 dvss.n70 dvss.n69 539.294
R4086 dvss.n2285 dvss.n70 539.294
R4087 dvss.n2285 dvss.n72 539.294
R4088 dvss.n73 dvss.n72 539.294
R4089 dvss.n2281 dvss.n73 539.294
R4090 dvss.n2281 dvss.n75 539.294
R4091 dvss.n76 dvss.n75 539.294
R4092 dvss.n1892 dvss.n76 539.294
R4093 dvss.n1892 dvss.n80 539.294
R4094 dvss.n81 dvss.n80 539.294
R4095 dvss.n1888 dvss.n81 539.294
R4096 dvss.n1888 dvss.n84 539.294
R4097 dvss.n85 dvss.n84 539.294
R4098 dvss.n203 dvss.n85 539.294
R4099 dvss.n203 dvss.n87 539.294
R4100 dvss.n88 dvss.n87 539.294
R4101 dvss.n199 dvss.n88 539.294
R4102 dvss.n199 dvss.n90 539.294
R4103 dvss.n91 dvss.n90 539.294
R4104 dvss.n195 dvss.n91 539.294
R4105 dvss.n195 dvss.n194 539.294
R4106 dvss.n194 dvss.n97 539.294
R4107 dvss.n98 dvss.n97 539.294
R4108 dvss.n189 dvss.n98 539.294
R4109 dvss.n189 dvss.n100 539.294
R4110 dvss.n101 dvss.n100 539.294
R4111 dvss.n185 dvss.n101 539.294
R4112 dvss.n185 dvss.n103 539.294
R4113 dvss.n104 dvss.n103 539.294
R4114 dvss.n181 dvss.n104 539.294
R4115 dvss.n181 dvss.n108 539.294
R4116 dvss.n109 dvss.n108 539.294
R4117 dvss.n171 dvss.n109 539.294
R4118 dvss.n171 dvss.n112 539.294
R4119 dvss.n113 dvss.n112 539.294
R4120 dvss.n174 dvss.n113 539.294
R4121 dvss.n174 dvss.n115 539.294
R4122 dvss.n116 dvss.n115 539.294
R4123 dvss.n118 dvss.n116 539.294
R4124 dvss.n3652 dvss.n118 539.294
R4125 dvss.n2277 dvss.n2276 503.457
R4126 dvss.n2278 dvss.n2277 503.457
R4127 dvss.n2290 dvss.n2289 503.457
R4128 dvss.n2288 dvss.n2287 503.457
R4129 dvss.n2287 dvss.n2286 503.457
R4130 dvss.n2286 dvss.n2284 503.457
R4131 dvss.n2229 dvss.n2228 503.457
R4132 dvss.n2230 dvss.n2229 503.457
R4133 dvss.n2234 dvss.n2231 503.457
R4134 dvss.n2236 dvss.n2235 503.457
R4135 dvss.n2238 dvss.n2236 503.457
R4136 dvss.n2239 dvss.n2238 503.457
R4137 dvss.n2240 dvss.n2239 503.457
R4138 dvss.n2242 dvss.n2240 503.457
R4139 dvss.n3649 dvss.n121 491.163
R4140 dvss.n2284 dvss.n2283 470.272
R4141 dvss.t62 dvss.n2278 445.769
R4142 dvss.t179 dvss.n2230 445.769
R4143 dvss.n3454 dvss.n3451 432.788
R4144 dvss.n3290 dvss.n250 432.788
R4145 dvss.n3173 dvss.n3172 432.788
R4146 dvss.n3056 dvss.n3055 432.788
R4147 dvss.n2943 dvss.n435 432.788
R4148 dvss.n1503 dvss.n1472 432.788
R4149 dvss.n1351 dvss.n544 432.788
R4150 dvss.n1091 dvss.n1090 432.788
R4151 dvss.n981 dvss.n751 432.788
R4152 dvss.n3450 dvss.t52 410.247
R4153 dvss.n3287 dvss.t26 410.247
R4154 dvss.n3171 dvss.t14 410.247
R4155 dvss.n3052 dvss.t4 410.247
R4156 dvss.n2930 dvss.t278 410.247
R4157 dvss.n1495 dvss.t372 410.247
R4158 dvss.n1338 dvss.t469 410.247
R4159 dvss.n1092 dvss.t246 410.247
R4160 dvss.n968 dvss.t72 410.247
R4161 dvss.t58 dvss.n3458 401.229
R4162 dvss.t32 dvss.n3309 401.229
R4163 dvss.n3190 dvss.t20 401.229
R4164 dvss.t10 dvss.n3077 401.229
R4165 dvss.n436 dvss.t274 401.229
R4166 dvss.t374 dvss.n1504 401.229
R4167 dvss.n545 dvss.t463 401.229
R4168 dvss.n646 dvss.t240 401.229
R4169 dvss.n982 dvss.t64 401.229
R4170 dvss.n3446 dvss.n3438 396.721
R4171 dvss.n269 dvss.n268 396.721
R4172 dvss.n333 dvss.n332 396.721
R4173 dvss.n391 dvss.n390 396.721
R4174 dvss.n2916 dvss.n2915 396.721
R4175 dvss.n1493 dvss.n1476 396.721
R4176 dvss.n1324 dvss.n1323 396.721
R4177 dvss.n1099 dvss.n1098 396.721
R4178 dvss.n959 dvss.n856 396.721
R4179 dvss.n2243 dvss.n2242 392.74
R4180 dvss.n2276 dvss.n2274 371.257
R4181 dvss.n2228 dvss.n2226 371.257
R4182 dvss.n3486 dvss.n121 358.591
R4183 dvss.n903 dvss.t310 349.909
R4184 dvss.n2220 dvss.n2219 344.817
R4185 dvss.n2226 dvss.n2225 344.817
R4186 dvss.n2244 dvss.n2243 344.817
R4187 dvss.n2265 dvss.n2264 344.817
R4188 dvss.n2268 dvss.n2267 344.817
R4189 dvss.n2274 dvss.n2273 344.817
R4190 dvss.n3470 dvss.n3420 332.075
R4191 dvss.n3486 dvss.n3485 332.075
R4192 dvss.n3337 dvss.n228 332.075
R4193 dvss.n3546 dvss.n207 332.075
R4194 dvss.n3224 dvss.n290 332.075
R4195 dvss.n3250 dvss.n3249 332.075
R4196 dvss.n3108 dvss.n354 332.075
R4197 dvss.n3134 dvss.n3133 332.075
R4198 dvss.n2989 dvss.n418 332.075
R4199 dvss.n3016 dvss.n3015 332.075
R4200 dvss.n1518 dvss.n1517 332.075
R4201 dvss.n2914 dvss.n449 332.075
R4202 dvss.n1397 dvss.n527 332.075
R4203 dvss.n1580 dvss.n506 332.075
R4204 dvss.n681 dvss.n680 332.075
R4205 dvss.n1322 dvss.n558 332.075
R4206 dvss.n1020 dvss.n733 332.075
R4207 dvss.n1107 dvss.n616 332.075
R4208 dvss.t135 dvss.n2263 308.899
R4209 dvss.n2289 dvss.t386 304.173
R4210 dvss.t432 dvss.n2234 304.173
R4211 dvss.n3458 dvss.t56 302.05
R4212 dvss.n3309 dvss.t30 302.05
R4213 dvss.n3190 dvss.t18 302.05
R4214 dvss.n3077 dvss.t8 302.05
R4215 dvss.t276 dvss.n436 302.05
R4216 dvss.n1504 dvss.t368 302.05
R4217 dvss.t465 dvss.n545 302.05
R4218 dvss.n646 dvss.t244 302.05
R4219 dvss.n982 dvss.t70 302.05
R4220 dvss.n3466 dvss.t300 297.485
R4221 dvss.n1887 dvss.t501 297.485
R4222 dvss.n3210 dvss.t224 297.485
R4223 dvss.n3094 dvss.t390 297.485
R4224 dvss.n1805 dvss.t189 297.485
R4225 dvss.n1514 dvss.t334 297.485
R4226 dvss.n1225 dvss.t408 297.485
R4227 dvss.n677 dvss.t424 297.485
R4228 dvss.n1005 dvss.t328 297.485
R4229 dvss.n2221 dvss.t534 294.531
R4230 dvss.n2269 dvss.t137 294.531
R4231 dvss.t54 dvss.n3450 293.034
R4232 dvss.n3287 dvss.t28 293.034
R4233 dvss.t16 dvss.n3171 293.034
R4234 dvss.n3052 dvss.t6 293.034
R4235 dvss.n2930 dvss.t280 293.034
R4236 dvss.n1495 dvss.t370 293.034
R4237 dvss.n1338 dvss.t467 293.034
R4238 dvss.n1092 dvss.t242 293.034
R4239 dvss.n968 dvss.t66 293.034
R4240 dvss.n3479 dvss.t302 283.649
R4241 dvss.n3343 dvss.t511 283.649
R4242 dvss.t226 dvss.n3228 283.649
R4243 dvss.t392 dvss.n3112 283.649
R4244 dvss.n2996 dvss.t185 283.649
R4245 dvss.n1525 dvss.t338 283.649
R4246 dvss.n1403 dvss.t400 283.649
R4247 dvss.n688 dvss.t420 283.649
R4248 dvss.n1026 dvss.t324 283.649
R4249 dvss.n3743 dvss.t347 282.327
R4250 dvss.n3749 dvss.t351 281.13
R4251 dvss.n3438 dvss.n207 276.731
R4252 dvss.n3250 dvss.n269 276.731
R4253 dvss.n3134 dvss.n333 276.731
R4254 dvss.n3016 dvss.n391 276.731
R4255 dvss.n2915 dvss.n2914 276.731
R4256 dvss.n1476 dvss.n506 276.731
R4257 dvss.n1323 dvss.n1322 276.731
R4258 dvss.n1099 dvss.n616 276.731
R4259 dvss.n2283 dvss.n2282 275.899
R4260 dvss.n2282 dvss.n2280 275.899
R4261 dvss.n2280 dvss.n2279 275.899
R4262 dvss.n2670 dvss.n2669 275.899
R4263 dvss.n204 dvss.n202 275.899
R4264 dvss.n202 dvss.n201 275.899
R4265 dvss.n201 dvss.n200 275.899
R4266 dvss.n200 dvss.n198 275.899
R4267 dvss.n198 dvss.n197 275.899
R4268 dvss.n196 dvss.n193 275.899
R4269 dvss.n192 dvss.n191 275.899
R4270 dvss.n191 dvss.n190 275.899
R4271 dvss.n190 dvss.n188 275.899
R4272 dvss.n188 dvss.n187 275.899
R4273 dvss.n187 dvss.n186 275.899
R4274 dvss.n186 dvss.n184 275.899
R4275 dvss.n184 dvss.n183 275.899
R4276 dvss.n180 dvss.n179 275.899
R4277 dvss.n175 dvss.n173 275.899
R4278 dvss.n173 dvss.n172 275.899
R4279 dvss.n172 dvss.n119 275.899
R4280 dvss.n3651 dvss.n119 275.899
R4281 dvss.n60 dvss.n9 270.307
R4282 dvss.n60 dvss.n10 270.307
R4283 dvss.n63 dvss.n9 270.307
R4284 dvss.n63 dvss.n10 270.307
R4285 dvss.t540 dvss.n2221 265.796
R4286 dvss.t145 dvss.n2269 265.796
R4287 dvss.t364 dvss.n3446 261.476
R4288 dvss.n268 dvss.t2 261.476
R4289 dvss.n332 dvss.t0 261.476
R4290 dvss.n390 dvss.t50 261.476
R4291 dvss.n2916 dvss.t84 261.476
R4292 dvss.t306 dvss.n1493 261.476
R4293 dvss.n1324 dvss.t248 261.476
R4294 dvss.n1098 dvss.t236 261.476
R4295 dvss.n959 dvss.t193 261.476
R4296 dvss.n2224 dvss.n2223 258.613
R4297 dvss.n2272 dvss.n2271 258.613
R4298 dvss.n3479 dvss.t298 255.976
R4299 dvss.n3343 dvss.t507 255.976
R4300 dvss.n3228 dvss.t234 255.976
R4301 dvss.n3112 dvss.t398 255.976
R4302 dvss.n2996 dvss.t181 255.976
R4303 dvss.n1525 dvss.t336 255.976
R4304 dvss.n1403 dvss.t402 255.976
R4305 dvss.n688 dvss.t418 255.976
R4306 dvss.n1026 dvss.t322 255.976
R4307 dvss.n3574 dvss.n3572 251.879
R4308 dvss.n3590 dvss.n3589 251.879
R4309 dvss.n3604 dvss.n147 251.879
R4310 dvss.n3606 dvss.n3605 251.879
R4311 dvss.n3606 dvss.n141 251.879
R4312 dvss.n3622 dvss.n141 251.879
R4313 dvss.n3624 dvss.n135 251.879
R4314 dvss.n3635 dvss.n135 251.879
R4315 dvss.n3638 dvss.n3637 251.879
R4316 dvss.n1851 dvss.n1850 251.879
R4317 dvss.n1855 dvss.n1854 251.879
R4318 dvss.n1858 dvss.n1857 251.879
R4319 dvss.n1861 dvss.n1860 251.879
R4320 dvss.n1862 dvss.n1861 251.879
R4321 dvss.n1863 dvss.n1862 251.879
R4322 dvss.n1868 dvss.n1867 251.879
R4323 dvss.n1870 dvss.n1868 251.879
R4324 dvss.n1873 dvss.n1872 251.879
R4325 dvss.n1881 dvss.n1880 251.879
R4326 dvss.n1885 dvss.n1884 251.879
R4327 dvss.n2673 dvss.n2672 251.879
R4328 dvss.n2676 dvss.n2675 251.879
R4329 dvss.n2677 dvss.n2676 251.879
R4330 dvss.n2679 dvss.n2677 251.879
R4331 dvss.n2681 dvss.n170 251.879
R4332 dvss.n3549 dvss.n170 251.879
R4333 dvss.n3570 dvss.n163 251.879
R4334 dvss.n1826 dvss.n1825 251.879
R4335 dvss.n1830 dvss.n1829 251.879
R4336 dvss.n1833 dvss.n1832 251.879
R4337 dvss.n1836 dvss.n1835 251.879
R4338 dvss.n1837 dvss.n1836 251.879
R4339 dvss.n1838 dvss.n1837 251.879
R4340 dvss.n1843 dvss.n1842 251.879
R4341 dvss.n1845 dvss.n1843 251.879
R4342 dvss.n1848 dvss.n1847 251.879
R4343 dvss.n1798 dvss.n1797 251.879
R4344 dvss.n1803 dvss.n1802 251.879
R4345 dvss.n1808 dvss.n1807 251.879
R4346 dvss.n1811 dvss.n1810 251.879
R4347 dvss.n1812 dvss.n1811 251.879
R4348 dvss.n1813 dvss.n1812 251.879
R4349 dvss.n1818 dvss.n1817 251.879
R4350 dvss.n1820 dvss.n1818 251.879
R4351 dvss.n1823 dvss.n1822 251.879
R4352 dvss.n1606 dvss.n1605 251.879
R4353 dvss.n1620 dvss.n486 251.879
R4354 dvss.n1623 dvss.n1622 251.879
R4355 dvss.n1636 dvss.n1635 251.879
R4356 dvss.n1638 dvss.n1636 251.879
R4357 dvss.n1638 dvss.n1637 251.879
R4358 dvss.n1652 dvss.n1651 251.879
R4359 dvss.n1652 dvss.n461 251.879
R4360 dvss.n2880 dvss.n462 251.879
R4361 dvss.n1218 dvss.n1217 251.879
R4362 dvss.n1223 dvss.n1222 251.879
R4363 dvss.n1228 dvss.n1227 251.879
R4364 dvss.n1231 dvss.n1230 251.879
R4365 dvss.n1232 dvss.n1231 251.879
R4366 dvss.n1233 dvss.n1232 251.879
R4367 dvss.n1238 dvss.n1237 251.879
R4368 dvss.n1238 dvss.n503 251.879
R4369 dvss.n1584 dvss.n1583 251.879
R4370 dvss.n1133 dvss.n1132 251.879
R4371 dvss.n1147 dvss.n596 251.879
R4372 dvss.n1150 dvss.n1149 251.879
R4373 dvss.n1163 dvss.n1162 251.879
R4374 dvss.n1165 dvss.n1163 251.879
R4375 dvss.n1165 dvss.n1164 251.879
R4376 dvss.n1179 dvss.n1178 251.879
R4377 dvss.n1179 dvss.n571 251.879
R4378 dvss.n1290 dvss.n572 251.879
R4379 dvss.n849 dvss.n765 251.879
R4380 dvss.n847 dvss.n773 251.879
R4381 dvss.n840 dvss.n839 251.879
R4382 dvss.n833 dvss.n806 251.879
R4383 dvss.n833 dvss.n832 251.879
R4384 dvss.n832 dvss.n831 251.879
R4385 dvss.n825 dvss.n824 251.879
R4386 dvss.n824 dvss.n613 251.879
R4387 dvss.n1111 dvss.n1110 251.879
R4388 dvss.n3482 dvss.n134 249.058
R4389 dvss.n3547 dvss.n205 249.058
R4390 dvss.n3227 dvss.n272 249.058
R4391 dvss.n3111 dvss.n336 249.058
R4392 dvss.n2995 dvss.n398 249.058
R4393 dvss.n2883 dvss.n2882 249.058
R4394 dvss.n1581 dvss.n504 249.058
R4395 dvss.n1293 dvss.n1292 249.058
R4396 dvss.n1108 dvss.n614 249.058
R4397 dvss.t487 dvss.n1893 247.16
R4398 dvss.n182 dvss.t99 247.16
R4399 dvss.t350 dvss 246.194
R4400 dvss.n1988 dvss.t313 245.276
R4401 dvss.n197 dvss.t109 244.286
R4402 dvss.n7 dvss.t428 236.149
R4403 dvss.n3572 dvss.n3571 230.888
R4404 dvss.n1850 dvss.n1849 230.888
R4405 dvss.n1880 dvss.n1879 230.888
R4406 dvss.n1825 dvss.n1824 230.888
R4407 dvss.n1797 dvss.n1796 230.888
R4408 dvss.n1605 dvss.n494 230.888
R4409 dvss.n1217 dvss.n1216 230.888
R4410 dvss.n1132 dvss.n604 230.888
R4411 dvss.n856 dvss.n765 230.888
R4412 dvss.n1134 dvss.t129 226.6
R4413 dvss.t485 dvss.n3573 226.6
R4414 dvss.n1853 dvss.t440 226.6
R4415 dvss.n1883 dvss.t522 226.6
R4416 dvss.n1828 dvss.t352 226.6
R4417 dvss.n1801 dvss.t289 226.6
R4418 dvss.n1607 dvss.t201 226.6
R4419 dvss.n1221 dvss.t220 226.6
R4420 dvss.t42 dvss.n848 226.6
R4421 dvss.n3591 dvss.t481 221.619
R4422 dvss.t446 dvss.n1856 221.619
R4423 dvss.t528 dvss.n1886 221.619
R4424 dvss.t358 dvss.n1831 221.619
R4425 dvss.t285 dvss.n1804 221.619
R4426 dvss.t203 dvss.n1621 221.619
R4427 dvss.t214 dvss.n1224 221.619
R4428 dvss.t133 dvss.n1148 221.619
R4429 dvss.n841 dvss.t44 221.619
R4430 dvss.n178 dvss.n177 220.345
R4431 dvss.n1891 dvss.n1890 220.345
R4432 dvss.n673 dvss.n645 217.097
R4433 dvss.n3460 dvss.n3459 217.097
R4434 dvss.n3311 dvss.n3310 217.097
R4435 dvss.n3195 dvss.n3194 217.097
R4436 dvss.n3079 dvss.n3078 217.097
R4437 dvss.n2963 dvss.n2962 217.097
R4438 dvss.n1505 dvss.n1470 217.097
R4439 dvss.n1371 dvss.n1370 217.097
R4440 dvss.n986 dvss.n748 217.097
R4441 dvss.n2263 dvss.n296 211.918
R4442 dvss.n3638 dvss.n120 209.899
R4443 dvss.n1879 dvss.n1873 209.899
R4444 dvss.n3571 dvss.n3570 209.899
R4445 dvss.n1849 dvss.n1848 209.899
R4446 dvss.n1824 dvss.n1823 209.899
R4447 dvss.n1796 dvss.n462 209.899
R4448 dvss.n1583 dvss.n494 209.899
R4449 dvss.n1216 dvss.n572 209.899
R4450 dvss.n1110 dvss.n604 209.899
R4451 dvss.n3747 dvss.n2 207.213
R4452 dvss.n24 dvss.n23 207.213
R4453 dvss.n28 dvss.n22 207.213
R4454 dvss.n31 dvss.n30 207.213
R4455 dvss.n37 dvss.n19 207.213
R4456 dvss.n40 dvss.n39 207.213
R4457 dvss.n17 dvss.n16 207.213
R4458 dvss.n51 dvss.n45 207.213
R4459 dvss.n3466 dvss.n146 204.089
R4460 dvss.n2671 dvss.n1887 204.089
R4461 dvss.n3210 dvss.n296 204.089
R4462 dvss.n3094 dvss.n360 204.089
R4463 dvss.n1806 dvss.n1805 204.089
R4464 dvss.n1514 dvss.n1513 204.089
R4465 dvss.n1226 dvss.n1225 204.089
R4466 dvss.n677 dvss.n676 204.089
R4467 dvss.n1005 dvss.n1004 204.089
R4468 dvss.n1893 dvss.t491 201.177
R4469 dvss.t95 dvss.n182 201.177
R4470 dvss.n1311 dvss.n557 200.215
R4471 dvss.n1488 dvss.n1487 200.215
R4472 dvss.n1489 dvss.n1488 200.215
R4473 dvss.n2900 dvss.n448 200.215
R4474 dvss.n2903 dvss.n448 200.215
R4475 dvss.n3035 dvss.n3034 200.215
R4476 dvss.n3036 dvss.n3035 200.215
R4477 dvss.n3138 dvss.n3137 200.215
R4478 dvss.n3139 dvss.n3138 200.215
R4479 dvss.n3254 dvss.n3253 200.215
R4480 dvss.n3255 dvss.n3254 200.215
R4481 dvss.n3437 dvss.n3436 200.215
R4482 dvss.n3437 dvss.n3432 200.215
R4483 dvss.n1101 dvss.n1100 200.215
R4484 dvss.n1100 dvss.n625 200.215
R4485 dvss.n1215 dvss.n1214 200.215
R4486 dvss.n1215 dvss.n1213 200.215
R4487 dvss.n1594 dvss.n1593 200.215
R4488 dvss.n1595 dvss.n1594 200.215
R4489 dvss.n1795 dvss.n1794 200.215
R4490 dvss.n1795 dvss.n1793 200.215
R4491 dvss.n1790 dvss.n1789 200.215
R4492 dvss.n1790 dvss.n1787 200.215
R4493 dvss.n1784 dvss.n1783 200.215
R4494 dvss.n1784 dvss.n1781 200.215
R4495 dvss.n1878 dvss.n1877 200.215
R4496 dvss.n1878 dvss.n1875 200.215
R4497 dvss.n3554 dvss.n162 200.215
R4498 dvss.n3557 dvss.n162 200.215
R4499 dvss.n1121 dvss.n1120 200.215
R4500 dvss.n1122 dvss.n1121 200.215
R4501 dvss.n1046 dvss.n717 200.215
R4502 dvss.n717 dvss.n716 200.215
R4503 dvss.n1307 dvss.n1306 200.215
R4504 dvss.n1306 dvss.n1305 200.215
R4505 dvss.n1480 dvss.n1479 200.215
R4506 dvss.n1481 dvss.n1480 200.215
R4507 dvss.n2896 dvss.n2895 200.215
R4508 dvss.n2895 dvss.n2894 200.215
R4509 dvss.n3023 dvss.n3022 200.215
R4510 dvss.n3024 dvss.n3023 200.215
R4511 dvss.n3148 dvss.n3147 200.215
R4512 dvss.n3149 dvss.n3148 200.215
R4513 dvss.n3264 dvss.n3263 200.215
R4514 dvss.n3265 dvss.n3264 200.215
R4515 dvss.n3442 dvss.n3441 200.215
R4516 dvss.n3443 dvss.n3442 200.215
R4517 dvss.n946 dvss.n863 200.215
R4518 dvss.n2666 dvss.n1895 200.215
R4519 dvss.n2666 dvss.n1896 200.215
R4520 dvss.n2666 dvss.n1897 200.215
R4521 dvss.n2666 dvss.n1898 200.215
R4522 dvss.n2666 dvss.n1899 200.215
R4523 dvss.n2666 dvss.n1900 200.215
R4524 dvss.n2666 dvss.n1901 200.215
R4525 dvss.n2666 dvss.n1902 200.215
R4526 dvss.n2666 dvss.n1903 200.215
R4527 dvss.n2666 dvss.n1904 200.215
R4528 dvss.n2666 dvss.n1905 200.215
R4529 dvss.n2666 dvss.n1906 200.215
R4530 dvss.n2666 dvss.n1907 200.215
R4531 dvss.n2666 dvss.n1908 200.215
R4532 dvss.n2666 dvss.n1909 200.215
R4533 dvss.n2666 dvss.n1910 200.215
R4534 dvss.n2666 dvss.n1911 200.215
R4535 dvss.n2666 dvss.n1912 200.215
R4536 dvss.n2666 dvss.n1913 200.215
R4537 dvss.n2666 dvss.n1914 200.215
R4538 dvss.n2666 dvss.n1915 200.215
R4539 dvss.n2666 dvss.n1916 200.215
R4540 dvss.n2666 dvss.n1917 200.215
R4541 dvss.n2666 dvss.n1918 200.215
R4542 dvss.n2666 dvss.n1919 200.215
R4543 dvss.n2666 dvss.n1920 200.215
R4544 dvss.n2666 dvss.n1921 200.215
R4545 dvss.n2666 dvss.n1922 200.215
R4546 dvss.n2666 dvss.n1923 200.215
R4547 dvss.n2666 dvss.n1924 200.215
R4548 dvss.n2666 dvss.n1925 200.215
R4549 dvss.n2666 dvss.n1926 200.215
R4550 dvss.n2666 dvss.n1927 200.215
R4551 dvss.n2666 dvss.n1928 200.215
R4552 dvss.n2666 dvss.n1929 200.215
R4553 dvss.n2666 dvss.n1930 200.215
R4554 dvss.n2666 dvss.n1931 200.215
R4555 dvss.n2666 dvss.n1932 200.215
R4556 dvss.n2666 dvss.n1933 200.215
R4557 dvss.n2666 dvss.n1934 200.215
R4558 dvss.n2666 dvss.n1935 200.215
R4559 dvss.n2666 dvss.n1936 200.215
R4560 dvss.n2666 dvss.n1937 200.215
R4561 dvss.n2666 dvss.n1938 200.215
R4562 dvss.n2666 dvss.n1939 200.215
R4563 dvss.n2666 dvss.n1940 200.215
R4564 dvss.n2666 dvss.n1941 200.215
R4565 dvss.n2666 dvss.n1942 200.215
R4566 dvss.n2666 dvss.n1943 200.215
R4567 dvss.n2666 dvss.n1944 200.215
R4568 dvss.n2666 dvss.n1945 200.215
R4569 dvss.n2666 dvss.n1946 200.215
R4570 dvss.n2666 dvss.n1947 200.215
R4571 dvss.n2666 dvss.n1948 200.215
R4572 dvss.n2666 dvss.n1949 200.215
R4573 dvss.n2666 dvss.n1950 200.215
R4574 dvss.n2666 dvss.n1951 200.215
R4575 dvss.n2666 dvss.n1952 200.215
R4576 dvss.n2666 dvss.n1953 200.215
R4577 dvss.n2666 dvss.n1954 200.215
R4578 dvss.n2666 dvss.n1955 200.215
R4579 dvss.n2666 dvss.n1956 200.215
R4580 dvss.n2666 dvss.n1957 200.215
R4581 dvss.n2666 dvss.n1958 200.215
R4582 dvss.n2666 dvss.n1959 200.215
R4583 dvss.n2666 dvss.n1960 200.215
R4584 dvss.n2666 dvss.n1961 200.215
R4585 dvss.n2666 dvss.n1962 200.215
R4586 dvss.n2666 dvss.n1963 200.215
R4587 dvss.t386 dvss.n2288 199.286
R4588 dvss.n2235 dvss.t432 199.286
R4589 dvss.n3636 dvss.n3635 188.91
R4590 dvss.n1871 dvss.n1870 188.91
R4591 dvss.n3549 dvss.n3548 188.91
R4592 dvss.n1846 dvss.n1845 188.91
R4593 dvss.n1821 dvss.n1820 188.91
R4594 dvss.n2881 dvss.n461 188.91
R4595 dvss.n1582 dvss.n503 188.91
R4596 dvss.n1291 dvss.n571 188.91
R4597 dvss.n1109 dvss.n613 188.91
R4598 dvss.t101 dvss.n176 188.212
R4599 dvss.t497 dvss.n1889 188.212
R4600 dvss.n1987 dvss.n1986 185
R4601 dvss.n946 dvss.n945 184.572
R4602 dvss.n1102 dvss.n1101 184.572
R4603 dvss.n628 dvss.n625 184.572
R4604 dvss.n1311 dvss.n1310 184.572
R4605 dvss.n1487 dvss.n1486 184.572
R4606 dvss.n1490 dvss.n1489 184.572
R4607 dvss.n2900 dvss.n452 184.572
R4608 dvss.n2903 dvss.n2902 184.572
R4609 dvss.n3034 dvss.n3033 184.572
R4610 dvss.n3037 dvss.n3036 184.572
R4611 dvss.n3137 dvss.n3136 184.572
R4612 dvss.n3139 dvss.n331 184.572
R4613 dvss.n3253 dvss.n3252 184.572
R4614 dvss.n3255 dvss.n267 184.572
R4615 dvss.n3436 dvss.n3435 184.572
R4616 dvss.n3432 dvss.n3431 184.572
R4617 dvss.n1312 dvss.n1311 184.572
R4618 dvss.n1487 dvss.n1485 184.572
R4619 dvss.n1489 dvss.n1484 184.572
R4620 dvss.n2901 dvss.n2900 184.572
R4621 dvss.n2904 dvss.n2903 184.572
R4622 dvss.n3034 dvss.n392 184.572
R4623 dvss.n3036 dvss.n389 184.572
R4624 dvss.n3137 dvss.n330 184.572
R4625 dvss.n3140 dvss.n3139 184.572
R4626 dvss.n3253 dvss.n266 184.572
R4627 dvss.n3256 dvss.n3255 184.572
R4628 dvss.n3436 dvss.n3434 184.572
R4629 dvss.n3433 dvss.n3432 184.572
R4630 dvss.n1101 dvss.n624 184.572
R4631 dvss.n1050 dvss.n625 184.572
R4632 dvss.n1120 dvss.n1119 184.572
R4633 dvss.n1123 dvss.n1122 184.572
R4634 dvss.n1214 dvss.n1184 184.572
R4635 dvss.n1213 dvss.n1212 184.572
R4636 dvss.n1593 dvss.n1592 184.572
R4637 dvss.n1596 dvss.n1595 184.572
R4638 dvss.n1794 dvss.n1657 184.572
R4639 dvss.n1793 dvss.n1792 184.572
R4640 dvss.n1789 dvss.n1788 184.572
R4641 dvss.n1787 dvss.n1690 184.572
R4642 dvss.n1783 dvss.n1782 184.572
R4643 dvss.n1781 dvss.n1721 184.572
R4644 dvss.n1877 dvss.n1876 184.572
R4645 dvss.n1875 dvss.n1752 184.572
R4646 dvss.n3554 dvss.n165 184.572
R4647 dvss.n3557 dvss.n3556 184.572
R4648 dvss.n3641 dvss.n3640 184.572
R4649 dvss.n1214 dvss.n1185 184.572
R4650 dvss.n1213 dvss.n1187 184.572
R4651 dvss.n1593 dvss.n498 184.572
R4652 dvss.n1595 dvss.n495 184.572
R4653 dvss.n1794 dvss.n1658 184.572
R4654 dvss.n1793 dvss.n1660 184.572
R4655 dvss.n1789 dvss.n1689 184.572
R4656 dvss.n1787 dvss.n1786 184.572
R4657 dvss.n1783 dvss.n1720 184.572
R4658 dvss.n1781 dvss.n1780 184.572
R4659 dvss.n1877 dvss.n1751 184.572
R4660 dvss.n1875 dvss.n1874 184.572
R4661 dvss.n3555 dvss.n3554 184.572
R4662 dvss.n3558 dvss.n3557 184.572
R4663 dvss.n1120 dvss.n608 184.572
R4664 dvss.n1122 dvss.n605 184.572
R4665 dvss.n1046 dvss.n1045 184.572
R4666 dvss.n716 dvss.n713 184.572
R4667 dvss.n1307 dvss.n1303 184.572
R4668 dvss.n1305 dvss.n555 184.572
R4669 dvss.n1479 dvss.n1478 184.572
R4670 dvss.n1482 dvss.n1481 184.572
R4671 dvss.n2896 dvss.n2892 184.572
R4672 dvss.n2894 dvss.n446 184.572
R4673 dvss.n3022 dvss.n3018 184.572
R4674 dvss.n3024 dvss.n3020 184.572
R4675 dvss.n3147 dvss.n3146 184.572
R4676 dvss.n3150 dvss.n3149 184.572
R4677 dvss.n3263 dvss.n3262 184.572
R4678 dvss.n3266 dvss.n3265 184.572
R4679 dvss.n3441 dvss.n3440 184.572
R4680 dvss.n3444 dvss.n3443 184.572
R4681 dvss.n1047 dvss.n1046 184.572
R4682 dvss.n716 dvss.n715 184.572
R4683 dvss.n1308 dvss.n1307 184.572
R4684 dvss.n1305 dvss.n1304 184.572
R4685 dvss.n1479 dvss.n1422 184.572
R4686 dvss.n1481 dvss.n1423 184.572
R4687 dvss.n2897 dvss.n2896 184.572
R4688 dvss.n2894 dvss.n2893 184.572
R4689 dvss.n3022 dvss.n3019 184.572
R4690 dvss.n3025 dvss.n3024 184.572
R4691 dvss.n3147 dvss.n324 184.572
R4692 dvss.n3149 dvss.n322 184.572
R4693 dvss.n3263 dvss.n260 184.572
R4694 dvss.n3265 dvss.n258 184.572
R4695 dvss.n3441 dvss.n3362 184.572
R4696 dvss.n3443 dvss.n3363 184.572
R4697 dvss.n860 dvss.n858 184.572
R4698 dvss.n947 dvss.n946 184.572
R4699 dvss.n855 dvss.n766 184.572
R4700 dvss.n1965 dvss.n1895 184.572
R4701 dvss.n1968 dvss.n1896 184.572
R4702 dvss.n1971 dvss.n1897 184.572
R4703 dvss.n1973 dvss.n1898 184.572
R4704 dvss.n1976 dvss.n1899 184.572
R4705 dvss.n1982 dvss.n1900 184.572
R4706 dvss.n1984 dvss.n1901 184.572
R4707 dvss.n1992 dvss.n1902 184.572
R4708 dvss.n1994 dvss.n1903 184.572
R4709 dvss.n1996 dvss.n1904 184.572
R4710 dvss.n2002 dvss.n1905 184.572
R4711 dvss.n2005 dvss.n1906 184.572
R4712 dvss.n2007 dvss.n1907 184.572
R4713 dvss.n2010 dvss.n1908 184.572
R4714 dvss.n2015 dvss.n1909 184.572
R4715 dvss.n2017 dvss.n1910 184.572
R4716 dvss.n2021 dvss.n1911 184.572
R4717 dvss.n2024 dvss.n1912 184.572
R4718 dvss.n2026 dvss.n1913 184.572
R4719 dvss.n2029 dvss.n1914 184.572
R4720 dvss.n2035 dvss.n1915 184.572
R4721 dvss.n2038 dvss.n1916 184.572
R4722 dvss.n2041 dvss.n1917 184.572
R4723 dvss.n2043 dvss.n1918 184.572
R4724 dvss.n2046 dvss.n1919 184.572
R4725 dvss.n2051 dvss.n1920 184.572
R4726 dvss.n2053 dvss.n1921 184.572
R4727 dvss.n2057 dvss.n1922 184.572
R4728 dvss.n2060 dvss.n1923 184.572
R4729 dvss.n2062 dvss.n1924 184.572
R4730 dvss.n2065 dvss.n1925 184.572
R4731 dvss.n2071 dvss.n1926 184.572
R4732 dvss.n2074 dvss.n1927 184.572
R4733 dvss.n2077 dvss.n1928 184.572
R4734 dvss.n2079 dvss.n1929 184.572
R4735 dvss.n2082 dvss.n1930 184.572
R4736 dvss.n2087 dvss.n1931 184.572
R4737 dvss.n2089 dvss.n1932 184.572
R4738 dvss.n2093 dvss.n1933 184.572
R4739 dvss.n2096 dvss.n1934 184.572
R4740 dvss.n2098 dvss.n1935 184.572
R4741 dvss.n2101 dvss.n1936 184.572
R4742 dvss.n2107 dvss.n1937 184.572
R4743 dvss.n2110 dvss.n1938 184.572
R4744 dvss.n2113 dvss.n1939 184.572
R4745 dvss.n2115 dvss.n1940 184.572
R4746 dvss.n2118 dvss.n1941 184.572
R4747 dvss.n2123 dvss.n1942 184.572
R4748 dvss.n2125 dvss.n1943 184.572
R4749 dvss.n2129 dvss.n1944 184.572
R4750 dvss.n2132 dvss.n1945 184.572
R4751 dvss.n2134 dvss.n1946 184.572
R4752 dvss.n2137 dvss.n1947 184.572
R4753 dvss.n2143 dvss.n1948 184.572
R4754 dvss.n2146 dvss.n1949 184.572
R4755 dvss.n2149 dvss.n1950 184.572
R4756 dvss.n2151 dvss.n1951 184.572
R4757 dvss.n2154 dvss.n1952 184.572
R4758 dvss.n2159 dvss.n1953 184.572
R4759 dvss.n2161 dvss.n1954 184.572
R4760 dvss.n2165 dvss.n1955 184.572
R4761 dvss.n2168 dvss.n1956 184.572
R4762 dvss.n2170 dvss.n1957 184.572
R4763 dvss.n2173 dvss.n1958 184.572
R4764 dvss.n2179 dvss.n1959 184.572
R4765 dvss.n2182 dvss.n1960 184.572
R4766 dvss.n2185 dvss.n1961 184.572
R4767 dvss.n2187 dvss.n1962 184.572
R4768 dvss.n2190 dvss.n1963 184.572
R4769 dvss.n1967 dvss.n1895 184.572
R4770 dvss.n1970 dvss.n1896 184.572
R4771 dvss.n1972 dvss.n1897 184.572
R4772 dvss.n1975 dvss.n1898 184.572
R4773 dvss.n1981 dvss.n1899 184.572
R4774 dvss.n1983 dvss.n1900 184.572
R4775 dvss.n1991 dvss.n1901 184.572
R4776 dvss.n1993 dvss.n1902 184.572
R4777 dvss.n1995 dvss.n1903 184.572
R4778 dvss.n2001 dvss.n1904 184.572
R4779 dvss.n2004 dvss.n1905 184.572
R4780 dvss.n2006 dvss.n1906 184.572
R4781 dvss.n2009 dvss.n1907 184.572
R4782 dvss.n2014 dvss.n1908 184.572
R4783 dvss.n2016 dvss.n1909 184.572
R4784 dvss.n2020 dvss.n1910 184.572
R4785 dvss.n2023 dvss.n1911 184.572
R4786 dvss.n2025 dvss.n1912 184.572
R4787 dvss.n2028 dvss.n1913 184.572
R4788 dvss.n2034 dvss.n1914 184.572
R4789 dvss.n2037 dvss.n1915 184.572
R4790 dvss.n2040 dvss.n1916 184.572
R4791 dvss.n2042 dvss.n1917 184.572
R4792 dvss.n2045 dvss.n1918 184.572
R4793 dvss.n2050 dvss.n1919 184.572
R4794 dvss.n2052 dvss.n1920 184.572
R4795 dvss.n2056 dvss.n1921 184.572
R4796 dvss.n2059 dvss.n1922 184.572
R4797 dvss.n2061 dvss.n1923 184.572
R4798 dvss.n2064 dvss.n1924 184.572
R4799 dvss.n2070 dvss.n1925 184.572
R4800 dvss.n2073 dvss.n1926 184.572
R4801 dvss.n2076 dvss.n1927 184.572
R4802 dvss.n2078 dvss.n1928 184.572
R4803 dvss.n2081 dvss.n1929 184.572
R4804 dvss.n2086 dvss.n1930 184.572
R4805 dvss.n2088 dvss.n1931 184.572
R4806 dvss.n2092 dvss.n1932 184.572
R4807 dvss.n2095 dvss.n1933 184.572
R4808 dvss.n2097 dvss.n1934 184.572
R4809 dvss.n2100 dvss.n1935 184.572
R4810 dvss.n2106 dvss.n1936 184.572
R4811 dvss.n2109 dvss.n1937 184.572
R4812 dvss.n2112 dvss.n1938 184.572
R4813 dvss.n2114 dvss.n1939 184.572
R4814 dvss.n2117 dvss.n1940 184.572
R4815 dvss.n2122 dvss.n1941 184.572
R4816 dvss.n2124 dvss.n1942 184.572
R4817 dvss.n2128 dvss.n1943 184.572
R4818 dvss.n2131 dvss.n1944 184.572
R4819 dvss.n2133 dvss.n1945 184.572
R4820 dvss.n2136 dvss.n1946 184.572
R4821 dvss.n2142 dvss.n1947 184.572
R4822 dvss.n2145 dvss.n1948 184.572
R4823 dvss.n2148 dvss.n1949 184.572
R4824 dvss.n2150 dvss.n1950 184.572
R4825 dvss.n2153 dvss.n1951 184.572
R4826 dvss.n2158 dvss.n1952 184.572
R4827 dvss.n2160 dvss.n1953 184.572
R4828 dvss.n2164 dvss.n1954 184.572
R4829 dvss.n2167 dvss.n1955 184.572
R4830 dvss.n2169 dvss.n1956 184.572
R4831 dvss.n2172 dvss.n1957 184.572
R4832 dvss.n2178 dvss.n1958 184.572
R4833 dvss.n2181 dvss.n1959 184.572
R4834 dvss.n2184 dvss.n1960 184.572
R4835 dvss.n2186 dvss.n1961 184.572
R4836 dvss.n2189 dvss.n1962 184.572
R4837 dvss.n2191 dvss.n1963 184.572
R4838 dvss.t538 dvss.n1894 179.593
R4839 dvss.t143 dvss.n2265 179.593
R4840 dvss.t294 dvss.n3470 172.957
R4841 dvss.n3337 dvss.t509 172.957
R4842 dvss.t232 dvss.n3224 172.957
R4843 dvss.t396 dvss.n3108 172.957
R4844 dvss.n2989 dvss.t187 172.957
R4845 dvss.n1518 dvss.t340 172.957
R4846 dvss.n1397 dvss.t406 172.957
R4847 dvss.n681 dvss.t422 172.957
R4848 dvss.n1020 dvss.t326 172.957
R4849 dvss.n3447 dvss.t364 171.311
R4850 dvss.n3286 dvss.t2 171.311
R4851 dvss.n3168 dvss.t0 171.311
R4852 dvss.n3051 dvss.t50 171.311
R4853 dvss.n2929 dvss.t84 171.311
R4854 dvss.n1494 dvss.t306 171.311
R4855 dvss.n1337 dvss.t248 171.311
R4856 dvss.n1061 dvss.t236 171.311
R4857 dvss.t193 dvss.n857 171.311
R4858 dvss.n1889 dvss.t493 169.85
R4859 dvss.n176 dvss.t97 169.85
R4860 dvss.n3471 dvss.t107 169.498
R4861 dvss.t451 dvss.n3340 169.498
R4862 dvss.t453 dvss.n3225 169.498
R4863 dvss.t412 dvss.n3109 169.498
R4864 dvss.t513 dvss.n2992 169.498
R4865 dvss.n1521 dvss.t318 169.498
R4866 dvss.t438 dvss.n1400 169.498
R4867 dvss.n684 dvss.t105 169.498
R4868 dvss.t436 dvss.n1023 169.498
R4869 dvss.n1148 dvss.t127 166.838
R4870 dvss.n3591 dvss.t479 166.838
R4871 dvss.n1856 dvss.t444 166.838
R4872 dvss.n1886 dvss.t526 166.838
R4873 dvss.n1831 dvss.t356 166.838
R4874 dvss.n1804 dvss.t287 166.838
R4875 dvss.n1621 dvss.t197 166.838
R4876 dvss.n1224 dvss.t216 166.838
R4877 dvss.n841 dvss.t40 166.838
R4878 dvss.n193 dvss.t456 166.689
R4879 dvss.n2219 dvss.t538 165.225
R4880 dvss.n2267 dvss.t143 165.225
R4881 dvss.n3478 dvss.t107 162.579
R4882 dvss.n3341 dvss.t451 162.579
R4883 dvss.n3229 dvss.t453 162.579
R4884 dvss.n3113 dvss.t412 162.579
R4885 dvss.n2993 dvss.t513 162.579
R4886 dvss.n1524 dvss.t318 162.579
R4887 dvss.n1401 dvss.t438 162.579
R4888 dvss.n687 dvss.t105 162.579
R4889 dvss.n1024 dvss.t436 162.579
R4890 dvss.n3524 dvss 161.882
R4891 dvss.n245 dvss 161.882
R4892 dvss.n310 dvss 161.882
R4893 dvss.n3062 dvss 161.882
R4894 dvss.n432 dvss 161.882
R4895 dvss.n1558 dvss 161.882
R4896 dvss.n541 dvss 161.882
R4897 dvss.n1070 dvss 161.882
R4898 dvss.n975 dvss 161.882
R4899 dvss.n3582 dvss 161.882
R4900 dvss.n1762 dvss 161.882
R4901 dvss.n1731 dvss 161.882
R4902 dvss.n1700 dvss 161.882
R4903 dvss.n1669 dvss 161.882
R4904 dvss.n1614 dvss 161.882
R4905 dvss.n1196 dvss 161.882
R4906 dvss.n1141 dvss 161.882
R4907 dvss.n791 dvss 161.882
R4908 dvss.n3573 dvss.t477 161.857
R4909 dvss.t442 dvss.n1853 161.857
R4910 dvss.t524 dvss.n1883 161.857
R4911 dvss.t354 dvss.n1828 161.857
R4912 dvss.t291 dvss.n1801 161.857
R4913 dvss.n1607 dvss.t199 161.857
R4914 dvss.t218 dvss.n1221 161.857
R4915 dvss.n1134 dvss.t125 161.857
R4916 dvss.n848 dvss.t36 161.857
R4917 dvss.n25 dvss.t178 161.47
R4918 dvss.n914 dvss.t262 160.064
R4919 dvss.t159 dvss.t177 155.49
R4920 dvss.t171 dvss.t159 155.49
R4921 dvss.t151 dvss.t171 155.49
R4922 dvss.t175 dvss.t151 155.49
R4923 dvss.t163 dvss.t175 155.49
R4924 dvss.t165 dvss.t163 155.49
R4925 dvss.t155 dvss.t165 155.49
R4926 dvss.t161 dvss.t155 155.49
R4927 dvss.t147 dvss.t161 155.49
R4928 dvss.t169 dvss.t147 155.49
R4929 dvss.t173 dvss.t149 155.49
R4930 dvss.t153 dvss.t173 155.49
R4931 dvss.t167 dvss.t153 155.49
R4932 dvss.t157 dvss.t167 155.49
R4933 dvss.t348 dvss.t350 155.49
R4934 dvss.t499 dvss.t348 155.49
R4935 dvss.t346 dvss.t499 155.49
R4936 dvss.t304 dvss.n3622 154.8
R4937 dvss.n1863 dvss.t228 154.8
R4938 dvss.t503 dvss.n2679 154.8
R4939 dvss.n1838 dvss.t394 154.8
R4940 dvss.n1813 dvss.t183 154.8
R4941 dvss.n1637 dvss.t332 154.8
R4942 dvss.n1233 dvss.t404 154.8
R4943 dvss.n1164 dvss.t416 154.8
R4944 dvss.n831 dvss.t320 154.8
R4945 dvss.n911 dvss.t476 154.305
R4946 dvss.n46 dvss.t158 152.838
R4947 dvss.n3464 dvss.t60 148.743
R4948 dvss.n3315 dvss.t34 148.743
R4949 dvss.t22 dvss.n304 148.743
R4950 dvss.t12 dvss.n368 148.743
R4951 dvss.n2967 dvss.t272 148.743
R4952 dvss.n1512 dvss.t366 148.743
R4953 dvss.n1375 dvss.t461 148.743
R4954 dvss.n675 dvss.t238 148.743
R4955 dvss.n1003 dvss.t68 148.743
R4956 dvss.n12 dvss.n10 146.25
R4957 dvss.n59 dvss.n12 146.25
R4958 dvss.n11 dvss.n9 146.25
R4959 dvss.n13 dvss.n11 146.25
R4960 dvss dvss.t157 144.385
R4961 dvss.n179 dvss.t93 143.697
R4962 dvss.n3451 dvss.t54 139.755
R4963 dvss.n3290 dvss.t28 139.755
R4964 dvss.n3173 dvss.t16 139.755
R4965 dvss.n3056 dvss.t6 139.755
R4966 dvss.t280 dvss.n435 139.755
R4967 dvss.t370 dvss.n1472 139.755
R4968 dvss.t467 dvss.n544 139.755
R4969 dvss.t242 dvss.n1091 139.755
R4970 dvss.t66 dvss.n751 139.755
R4971 dvss.n1978 dvss.t311 139.52
R4972 dvss.t483 dvss.n3604 139.059
R4973 dvss.t448 dvss.n1858 139.059
R4974 dvss.t530 dvss.n2673 139.059
R4975 dvss.t360 dvss.n1833 139.059
R4976 dvss.t283 dvss.n1808 139.059
R4977 dvss.n1622 dvss.t195 139.059
R4978 dvss.t222 dvss.n1228 139.059
R4979 dvss.n1149 dvss.t131 139.059
R4980 dvss.n839 dvss.t38 139.059
R4981 dvss dvss.t346 138.831
R4982 dvss.n914 dvss.t260 137.442
R4983 dvss.n915 dvss.t258 137.442
R4984 dvss.n3460 dvss.t60 134.488
R4985 dvss.n3311 dvss.t34 134.488
R4986 dvss.n3195 dvss.t22 134.488
R4987 dvss.n3079 dvss.t12 134.488
R4988 dvss.n2963 dvss.t272 134.488
R4989 dvss.n1470 dvss.t366 134.488
R4990 dvss.n1371 dvss.t461 134.488
R4991 dvss.t238 dvss.n673 134.488
R4992 dvss.n986 dvss.t68 134.488
R4993 dvss.n3454 dvss.t56 130.738
R4994 dvss.n250 dvss.t30 130.738
R4995 dvss.n3172 dvss.t18 130.738
R4996 dvss.n3055 dvss.t8 130.738
R4997 dvss.n2943 dvss.t276 130.738
R4998 dvss.t368 dvss.n1503 130.738
R4999 dvss.n1351 dvss.t465 130.738
R5000 dvss.n1090 dvss.t244 130.738
R5001 dvss.t70 dvss.n981 130.738
R5002 dvss.t205 dvss.n3623 128.564
R5003 dvss.t376 dvss.n1866 128.564
R5004 dvss.t382 dvss.n2680 128.564
R5005 dvss.t378 dvss.n1841 128.564
R5006 dvss.t24 dvss.n1816 128.564
R5007 dvss.t362 dvss.n1650 128.564
R5008 dvss.t414 dvss.n1236 128.564
R5009 dvss.t250 dvss.n1177 128.564
R5010 dvss.t473 dvss.n823 128.564
R5011 dvss.n3471 dvss.t103 127.987
R5012 dvss.n3340 dvss.t489 127.987
R5013 dvss.n3225 dvss.t139 127.987
R5014 dvss.n3109 dvss.t536 127.987
R5015 dvss.n2992 dvss.t208 127.987
R5016 dvss.n1521 dvss.t263 127.987
R5017 dvss.n1400 dvss.t517 127.987
R5018 dvss.n684 dvss.t86 127.987
R5019 dvss.n1023 dvss.t76 127.987
R5020 dvss.t95 dvss.n146 125.389
R5021 dvss.n2671 dvss.t491 125.389
R5022 dvss.n900 dvss.n876 124.787
R5023 dvss.n894 dvss.n876 124.787
R5024 dvss.n894 dvss.n893 124.787
R5025 dvss.n893 dvss.n892 124.787
R5026 dvss.n892 dvss.n882 124.787
R5027 dvss.n882 dvss.n875 124.787
R5028 dvss.n906 dvss.n875 124.787
R5029 dvss.n923 dvss.n922 124.787
R5030 dvss.n925 dvss.n923 124.787
R5031 dvss.n942 dvss.n941 124.787
R5032 dvss.n943 dvss.n942 124.787
R5033 dvss.n2669 dvss.n2668 123.579
R5034 dvss.n3624 dvss.t205 123.316
R5035 dvss.n1867 dvss.t376 123.316
R5036 dvss.n2681 dvss.t382 123.316
R5037 dvss.n1842 dvss.t378 123.316
R5038 dvss.n1817 dvss.t24 123.316
R5039 dvss.n1651 dvss.t362 123.316
R5040 dvss.n1237 dvss.t414 123.316
R5041 dvss.n1178 dvss.t250 123.316
R5042 dvss.n825 dvss.t473 123.316
R5043 dvss.n924 dvss.t255 120.886
R5044 dvss.n922 dvss.t475 116.987
R5045 dvss.n3661 dvss.t98 116.939
R5046 dvss.n3708 dvss.t494 116.939
R5047 dvss.n2310 dvss.t146 116.939
R5048 dvss.n2357 dvss.t541 116.939
R5049 dvss.n2404 dvss.t207 116.939
R5050 dvss.n2451 dvss.t266 116.939
R5051 dvss.n2498 dvss.t516 116.939
R5052 dvss.n2545 dvss.t88 116.939
R5053 dvss.n2592 dvss.t79 116.939
R5054 dvss.n3496 dvss.t299 116.939
R5055 dvss.n3354 dvss.t508 116.939
R5056 dvss.n3240 dvss.t235 116.939
R5057 dvss.n3124 dvss.t399 116.939
R5058 dvss.n3007 dvss.t182 116.939
R5059 dvss.n2888 dvss.t337 116.939
R5060 dvss.n1414 dvss.t403 116.939
R5061 dvss.n1298 dvss.t419 116.939
R5062 dvss.n1038 dvss.t323 116.939
R5063 dvss.n3515 dvss.t61 116.938
R5064 dvss.n3320 dvss.t35 116.938
R5065 dvss.n3204 dvss.t23 116.938
R5066 dvss.n3088 dvss.t13 116.938
R5067 dvss.n2972 dvss.t273 116.938
R5068 dvss.n1549 dvss.t367 116.938
R5069 dvss.n1380 dvss.t462 116.938
R5070 dvss.n1078 dvss.t239 116.938
R5071 dvss.n997 dvss.t69 116.938
R5072 dvss.n3599 dvss.t484 116.938
R5073 dvss.n2697 dvss.t531 116.938
R5074 dvss.n2747 dvss.t449 116.938
R5075 dvss.n2797 dvss.t361 116.938
R5076 dvss.n2847 dvss.t284 116.938
R5077 dvss.n1630 dvss.t196 116.938
R5078 dvss.n1257 dvss.t223 116.938
R5079 dvss.n1157 dvss.t132 116.938
R5080 dvss.n801 dvss.t39 116.938
R5081 dvss.n1004 dvss.t78 116.547
R5082 dvss.n1226 dvss.t78 116.547
R5083 dvss.n1806 dvss.t78 116.547
R5084 dvss.n1513 dvss.t78 116.547
R5085 dvss.n676 dvss.t78 116.547
R5086 dvss dvss.n3398 113.316
R5087 dvss dvss.n3328 113.316
R5088 dvss dvss.n3217 113.316
R5089 dvss dvss.n3101 113.316
R5090 dvss dvss.n2980 113.316
R5091 dvss dvss.n1461 113.316
R5092 dvss dvss.n1388 113.316
R5093 dvss dvss.n663 113.316
R5094 dvss dvss.n1011 113.316
R5095 dvss dvss.n3612 113.316
R5096 dvss dvss.n1773 113.316
R5097 dvss dvss.n1742 113.316
R5098 dvss dvss.n1711 113.316
R5099 dvss dvss.n1680 113.316
R5100 dvss dvss.n471 113.316
R5101 dvss dvss.n1207 113.316
R5102 dvss dvss.n581 113.316
R5103 dvss dvss.n812 113.316
R5104 dvss.n3605 dvss.t483 112.822
R5105 dvss.n1860 dvss.t448 112.822
R5106 dvss.n2675 dvss.t530 112.822
R5107 dvss.n1835 dvss.t360 112.822
R5108 dvss.n1810 dvss.t283 112.822
R5109 dvss.n1635 dvss.t195 112.822
R5110 dvss.n1230 dvss.t222 112.822
R5111 dvss.n1162 dvss.t131 112.822
R5112 dvss.n806 dvss.t38 112.822
R5113 dvss.t456 dvss.n192 109.21
R5114 dvss.n935 dvss.n933 105.862
R5115 dvss.t495 dvss.n1891 105.582
R5116 dvss.t93 dvss.n178 105.582
R5117 dvss.t149 dvss.n57 99.9584
R5118 dvss.n3623 dvss.t304 97.0786
R5119 dvss.n1866 dvss.t228 97.0786
R5120 dvss.n2680 dvss.t503 97.0786
R5121 dvss.n1841 dvss.t394 97.0786
R5122 dvss.n1816 dvss.t183 97.0786
R5123 dvss.n1650 dvss.t332 97.0786
R5124 dvss.n1236 dvss.t404 97.0786
R5125 dvss.n1177 dvss.t416 97.0786
R5126 dvss.n823 dvss.t320 97.0786
R5127 dvss.n2244 dvss.t141 93.3883
R5128 dvss.t316 dvss.n856 92.29
R5129 dvss.n94 dvss.n93 90.0716
R5130 dvss.n2294 dvss.n2293 90.0716
R5131 dvss.n2208 dvss.n2207 90.0716
R5132 dvss.n2176 dvss.n2175 90.0716
R5133 dvss.n2140 dvss.n2139 90.0716
R5134 dvss.n2104 dvss.n2103 90.0716
R5135 dvss.n2068 dvss.n2067 90.0716
R5136 dvss.n2032 dvss.n2031 90.0716
R5137 dvss.n1999 dvss.n1998 90.0716
R5138 dvss.n1980 dvss.n1979 90.0716
R5139 dvss.n3368 dvss.n3367 90.0716
R5140 dvss.n3271 dvss.n3270 90.0716
R5141 dvss.n3156 dvss.n3155 90.0716
R5142 dvss.n3042 dvss.n3041 90.0716
R5143 dvss.n2923 dvss.n2922 90.0716
R5144 dvss.n1428 dvss.n1427 90.0716
R5145 dvss.n1331 dvss.n1330 90.0716
R5146 dvss.n1054 dvss.n1053 90.0716
R5147 dvss.n951 dvss.n950 90.0716
R5148 dvss.n3464 dvss.t296 89.9376
R5149 dvss.n3315 dvss.t505 89.9376
R5150 dvss.n304 dvss.t230 89.9376
R5151 dvss.n368 dvss.t388 89.9376
R5152 dvss.n2967 dvss.t191 89.9376
R5153 dvss.t342 dvss.n1512 89.9376
R5154 dvss.n1375 dvss.t410 89.9376
R5155 dvss.t426 dvss.n675 89.9376
R5156 dvss.t330 dvss.n1003 89.9376
R5157 dvss.n2225 dvss.n2224 86.2046
R5158 dvss.n2273 dvss.n2272 86.2046
R5159 dvss.n66 dvss.t112 84.171
R5160 dvss.n3485 dvss.n134 83.0194
R5161 dvss.n3547 dvss.n3546 83.0194
R5162 dvss.n3249 dvss.n272 83.0194
R5163 dvss.n3133 dvss.n336 83.0194
R5164 dvss.n3015 dvss.n398 83.0194
R5165 dvss.n2882 dvss.n449 83.0194
R5166 dvss.n1581 dvss.n1580 83.0194
R5167 dvss.n1292 dvss.n558 83.0194
R5168 dvss.n1108 dvss.n1107 83.0194
R5169 dvss.t257 dvss.n924 81.8912
R5170 dvss.n3589 dvss.t477 81.3362
R5171 dvss.n1854 dvss.t442 81.3362
R5172 dvss.n1884 dvss.t524 81.3362
R5173 dvss.n1829 dvss.t354 81.3362
R5174 dvss.n1802 dvss.t291 81.3362
R5175 dvss.n486 dvss.t199 81.3362
R5176 dvss.n1222 dvss.t218 81.3362
R5177 dvss.n596 dvss.t125 81.3362
R5178 dvss.t36 dvss.n847 81.3362
R5179 dvss.n2223 dvss.t540 79.0209
R5180 dvss.n2271 dvss.t145 79.0209
R5181 dvss.n901 dvss.n360 76.8976
R5182 dvss.n3678 dvss.n106 76.7239
R5183 dvss.n3661 dvss.n106 76.7239
R5184 dvss.n3725 dvss.n78 76.7239
R5185 dvss.n3708 dvss.n78 76.7239
R5186 dvss.n2327 dvss.n2247 76.7239
R5187 dvss.n2310 dvss.n2247 76.7239
R5188 dvss.n2374 dvss.n2193 76.7239
R5189 dvss.n2357 dvss.n2193 76.7239
R5190 dvss.n2421 dvss.n2156 76.7239
R5191 dvss.n2404 dvss.n2156 76.7239
R5192 dvss.n2468 dvss.n2120 76.7239
R5193 dvss.n2451 dvss.n2120 76.7239
R5194 dvss.n2515 dvss.n2084 76.7239
R5195 dvss.n2498 dvss.n2084 76.7239
R5196 dvss.n2562 dvss.n2048 76.7239
R5197 dvss.n2545 dvss.n2048 76.7239
R5198 dvss.n2609 dvss.n2012 76.7239
R5199 dvss.n2592 dvss.n2012 76.7239
R5200 dvss.n3497 dvss.n3403 76.7239
R5201 dvss.n3497 dvss.n3496 76.7239
R5202 dvss.n3353 dvss.n216 76.7239
R5203 dvss.n3354 dvss.n3353 76.7239
R5204 dvss.n3239 dvss.n279 76.7239
R5205 dvss.n3240 dvss.n3239 76.7239
R5206 dvss.n3123 dvss.n343 76.7239
R5207 dvss.n3124 dvss.n3123 76.7239
R5208 dvss.n3006 dvss.n406 76.7239
R5209 dvss.n3007 dvss.n3006 76.7239
R5210 dvss.n1456 dvss.n457 76.7239
R5211 dvss.n2888 dvss.n457 76.7239
R5212 dvss.n1413 dvss.n515 76.7239
R5213 dvss.n1414 dvss.n1413 76.7239
R5214 dvss.n658 dvss.n567 76.7239
R5215 dvss.n1298 dvss.n567 76.7239
R5216 dvss.n1036 dvss.n721 76.7239
R5217 dvss.n1038 dvss.n1036 76.7239
R5218 dvss.n906 dvss.n905 76.6918
R5219 dvss.n3482 dvss.t298 76.1011
R5220 dvss.t507 dvss.n205 76.1011
R5221 dvss.t234 dvss.n3227 76.1011
R5222 dvss.t398 dvss.n3111 76.1011
R5223 dvss.t181 dvss.n2995 76.1011
R5224 dvss.n2883 dvss.t336 76.1011
R5225 dvss.t402 dvss.n504 76.1011
R5226 dvss.n1293 dvss.t418 76.1011
R5227 dvss.t322 dvss.n614 76.1011
R5228 dvss.t479 dvss.n3590 76.0887
R5229 dvss.t444 dvss.n1855 76.0887
R5230 dvss.t526 dvss.n1885 76.0887
R5231 dvss.t356 dvss.n1830 76.0887
R5232 dvss.t287 dvss.n1803 76.0887
R5233 dvss.t197 dvss.n1620 76.0887
R5234 dvss.t216 dvss.n1223 76.0887
R5235 dvss.t127 dvss.n1147 76.0887
R5236 dvss.n773 dvss.t40 76.0887
R5237 dvss.n2279 dvss.t491 74.7229
R5238 dvss.n183 dvss.t95 74.7229
R5239 dvss dvss.n3524 73.0358
R5240 dvss.n3514 dvss 73.0358
R5241 dvss dvss.n245 73.0358
R5242 dvss dvss.n3299 73.0358
R5243 dvss dvss.n310 73.0358
R5244 dvss dvss.n3184 73.0358
R5245 dvss.n3062 dvss 73.0358
R5246 dvss dvss.n3064 73.0358
R5247 dvss dvss.n432 73.0358
R5248 dvss dvss.n2951 73.0358
R5249 dvss dvss.n1558 73.0358
R5250 dvss.n1548 dvss 73.0358
R5251 dvss dvss.n541 73.0358
R5252 dvss dvss.n1359 73.0358
R5253 dvss.n1070 dvss 73.0358
R5254 dvss.n1077 dvss 73.0358
R5255 dvss.n975 dvss 73.0358
R5256 dvss.n996 dvss 73.0358
R5257 dvss.n3582 dvss 73.0358
R5258 dvss.n3598 dvss 73.0358
R5259 dvss.n1762 dvss 73.0358
R5260 dvss.n2696 dvss 73.0358
R5261 dvss.n1731 dvss 73.0358
R5262 dvss.n2746 dvss 73.0358
R5263 dvss.n1700 dvss 73.0358
R5264 dvss.n2796 dvss 73.0358
R5265 dvss.n1669 dvss 73.0358
R5266 dvss.n2846 dvss 73.0358
R5267 dvss.n1614 dvss 73.0358
R5268 dvss.n1629 dvss 73.0358
R5269 dvss.n1196 dvss 73.0358
R5270 dvss.n1256 dvss 73.0358
R5271 dvss.n1141 dvss 73.0358
R5272 dvss.n1156 dvss 73.0358
R5273 dvss.n791 dvss 73.0358
R5274 dvss.n799 dvss 73.0358
R5275 dvss.n8 dvss.n6 66.771
R5276 dvss.n65 dvss.n5 66.771
R5277 dvss.n859 dvss.t459 65.1619
R5278 dvss.n3439 dvss.t252 64.6673
R5279 dvss.n259 dvss.t471 64.6673
R5280 dvss.n323 dvss.t542 64.6673
R5281 dvss.n3021 dvss.t46 64.6673
R5282 dvss.n447 dvss.t123 64.6673
R5283 dvss.n1477 dvss.t270 64.6673
R5284 dvss.n556 dvss.t121 64.6673
R5285 dvss.n626 dvss.t48 64.6673
R5286 dvss.t493 dvss.n204 63.2272
R5287 dvss.t97 dvss.n175 63.2272
R5288 dvss.n3637 dvss.n3636 62.9701
R5289 dvss.n1872 dvss.n1871 62.9701
R5290 dvss.n3548 dvss.n163 62.9701
R5291 dvss.n1847 dvss.n1846 62.9701
R5292 dvss.n1822 dvss.n1821 62.9701
R5293 dvss.n2881 dvss.n2880 62.9701
R5294 dvss.n1584 dvss.n1582 62.9701
R5295 dvss.n1291 dvss.n1290 62.9701
R5296 dvss.n1111 dvss.n1109 62.9701
R5297 dvss.n2666 dvss.t74 58.6242
R5298 dvss.n2290 dvss.t62 57.6882
R5299 dvss.n2231 dvss.t179 57.6882
R5300 dvss.n3678 dvss.n3677 57.0829
R5301 dvss.n3670 dvss.n3669 57.0829
R5302 dvss.n3725 dvss.n3724 57.0829
R5303 dvss.n3717 dvss.n3716 57.0829
R5304 dvss.n2327 dvss.n2326 57.0829
R5305 dvss.n2319 dvss.n2318 57.0829
R5306 dvss.n2374 dvss.n2373 57.0829
R5307 dvss.n2366 dvss.n2365 57.0829
R5308 dvss.n2421 dvss.n2420 57.0829
R5309 dvss.n2413 dvss.n2412 57.0829
R5310 dvss.n2468 dvss.n2467 57.0829
R5311 dvss.n2460 dvss.n2459 57.0829
R5312 dvss.n2515 dvss.n2514 57.0829
R5313 dvss.n2507 dvss.n2506 57.0829
R5314 dvss.n2562 dvss.n2561 57.0829
R5315 dvss.n2554 dvss.n2553 57.0829
R5316 dvss.n2609 dvss.n2608 57.0829
R5317 dvss.n2601 dvss.n2600 57.0829
R5318 dvss.n3403 dvss.n3402 57.0829
R5319 dvss.n3500 dvss.n3498 57.0829
R5320 dvss.n216 dvss.n215 57.0829
R5321 dvss.n3352 dvss.n218 57.0829
R5322 dvss.n279 dvss.n278 57.0829
R5323 dvss.n3238 dvss.n281 57.0829
R5324 dvss.n343 dvss.n342 57.0829
R5325 dvss.n3122 dvss.n345 57.0829
R5326 dvss.n406 dvss.n405 57.0829
R5327 dvss.n3005 dvss.n408 57.0829
R5328 dvss.n1456 dvss.n1455 57.0829
R5329 dvss.n1534 dvss.n1532 57.0829
R5330 dvss.n515 dvss.n514 57.0829
R5331 dvss.n1412 dvss.n517 57.0829
R5332 dvss.n658 dvss.n657 57.0829
R5333 dvss.n697 dvss.n695 57.0829
R5334 dvss.n721 dvss.n720 57.0829
R5335 dvss.n1035 dvss.n723 57.0829
R5336 dvss.n57 dvss.t169 55.5327
R5337 dvss.t534 dvss.n2220 50.2862
R5338 dvss.t137 dvss.n2268 50.2862
R5339 dvss.t302 dvss.n3478 48.4282
R5340 dvss.t511 dvss.n3341 48.4282
R5341 dvss.n3229 dvss.t226 48.4282
R5342 dvss.n3113 dvss.t392 48.4282
R5343 dvss.t185 dvss.n2993 48.4282
R5344 dvss.t338 dvss.n1524 48.4282
R5345 dvss.t400 dvss.n1401 48.4282
R5346 dvss.t420 dvss.n687 48.4282
R5347 dvss.t324 dvss.n1024 48.4282
R5348 dvss.n905 dvss.n904 48.095
R5349 dvss.n3378 dvss.n3377 46.2505
R5350 dvss.n3380 dvss.n3379 46.2505
R5351 dvss.n3281 dvss.n3277 46.2505
R5352 dvss.n3298 dvss.n3297 46.2505
R5353 dvss.n3163 dvss.n3159 46.2505
R5354 dvss.n3183 dvss.n3182 46.2505
R5355 dvss.n377 dvss.n376 46.2505
R5356 dvss.n3068 dvss.n3063 46.2505
R5357 dvss.n2936 dvss.n2935 46.2505
R5358 dvss.n2950 dvss.n2949 46.2505
R5359 dvss.n1438 dvss.n1437 46.2505
R5360 dvss.n1440 dvss.n1439 46.2505
R5361 dvss.n1344 dvss.n1343 46.2505
R5362 dvss.n1358 dvss.n1357 46.2505
R5363 dvss.n711 dvss.n710 46.2505
R5364 dvss.n1074 dvss.n1073 46.2505
R5365 dvss.n757 dvss.n756 46.2505
R5366 dvss.n744 dvss.n743 46.2505
R5367 dvss.n159 dvss.n158 46.2505
R5368 dvss.n153 dvss.n152 46.2505
R5369 dvss.n2714 dvss.n1757 46.2505
R5370 dvss.n2705 dvss.n1763 46.2505
R5371 dvss.n2764 dvss.n1726 46.2505
R5372 dvss.n2755 dvss.n1732 46.2505
R5373 dvss.n2814 dvss.n1695 46.2505
R5374 dvss.n2805 dvss.n1701 46.2505
R5375 dvss.n2864 dvss.n1663 46.2505
R5376 dvss.n2855 dvss.n1670 46.2505
R5377 dvss.n491 dvss.n490 46.2505
R5378 dvss.n482 dvss.n481 46.2505
R5379 dvss.n1274 dvss.n1190 46.2505
R5380 dvss.n1265 dvss.n1197 46.2505
R5381 dvss.n601 dvss.n600 46.2505
R5382 dvss.n592 dvss.n591 46.2505
R5383 dvss.n785 dvss.n784 46.2505
R5384 dvss.n795 dvss.n794 46.2505
R5385 dvss.n63 dvss.n62 45.0005
R5386 dvss.n62 dvss.t344 45.0005
R5387 dvss.n61 dvss.n60 45.0005
R5388 dvss.t344 dvss.n61 45.0005
R5389 dvss.n57 dvss.n56 45.0005
R5390 dvss.n3514 dvss 44.424
R5391 dvss.n3299 dvss 44.424
R5392 dvss.n3184 dvss 44.424
R5393 dvss.n3064 dvss 44.424
R5394 dvss.n2951 dvss 44.424
R5395 dvss.n1548 dvss 44.424
R5396 dvss.n1359 dvss 44.424
R5397 dvss.n1077 dvss 44.424
R5398 dvss.n996 dvss 44.424
R5399 dvss.n3598 dvss 44.424
R5400 dvss.n2696 dvss 44.424
R5401 dvss.n2746 dvss 44.424
R5402 dvss.n2796 dvss 44.424
R5403 dvss.n2846 dvss 44.424
R5404 dvss.n1629 dvss 44.424
R5405 dvss.n1256 dvss 44.424
R5406 dvss.n1156 dvss 44.424
R5407 dvss.n799 dvss 44.424
R5408 dvss.t313 dvss.n1987 43.2419
R5409 dvss.n925 dvss.t257 42.8956
R5410 dvss.t141 dvss.n296 39.5107
R5411 dvss.t296 dvss.n146 38.0508
R5412 dvss.n2671 dvss.t505 38.0508
R5413 dvss.t230 dvss.n296 38.0508
R5414 dvss.t388 dvss.n360 38.0508
R5415 dvss.n1806 dvss.t191 38.0508
R5416 dvss.n1513 dvss.t342 38.0508
R5417 dvss.n1226 dvss.t410 38.0508
R5418 dvss.n676 dvss.t426 38.0508
R5419 dvss.n1004 dvss.t330 38.0508
R5420 dvss.n933 dvss.t317 37.7206
R5421 dvss.n898 dvss.n897 36.1417
R5422 dvss.n897 dvss.n896 36.1417
R5423 dvss.n896 dvss.n880 36.1417
R5424 dvss.n890 dvss.n880 36.1417
R5425 dvss.n890 dvss.n889 36.1417
R5426 dvss.n889 dvss.n873 36.1417
R5427 dvss.n908 dvss.n873 36.1417
R5428 dvss.n908 dvss.n872 36.1417
R5429 dvss.n920 dvss.n872 36.1417
R5430 dvss.n920 dvss.n869 36.1417
R5431 dvss.n927 dvss.n869 36.1417
R5432 dvss.n927 dvss.n867 36.1417
R5433 dvss.n939 dvss.n867 36.1417
R5434 dvss.n939 dvss.n938 36.1417
R5435 dvss.n938 dvss.n865 36.1417
R5436 dvss.n865 dvss.n862 36.1417
R5437 dvss.n948 dvss.n862 36.1417
R5438 dvss.n948 dvss.n762 36.1417
R5439 dvss.n961 dvss.n762 36.1417
R5440 dvss.n962 dvss.n961 36.1417
R5441 dvss.n962 dvss.n758 36.1417
R5442 dvss.n971 dvss.n758 36.1417
R5443 dvss.n971 dvss.n754 36.1417
R5444 dvss.n754 dvss.n750 36.1417
R5445 dvss.n750 dvss.n745 36.1417
R5446 dvss.n985 dvss.n745 36.1417
R5447 dvss.n985 dvss.n736 36.1417
R5448 dvss.n1007 dvss.n736 36.1417
R5449 dvss.n1008 dvss.n1007 36.1417
R5450 dvss.n1008 dvss.n732 36.1417
R5451 dvss.n732 dvss.n724 36.1417
R5452 dvss.n729 dvss.n724 36.1417
R5453 dvss.n1028 dvss.n729 36.1417
R5454 dvss.n1028 dvss.n619 36.1417
R5455 dvss.n1105 dvss.n619 36.1417
R5456 dvss.n1105 dvss.n1104 36.1417
R5457 dvss.n1104 dvss.n1103 36.1417
R5458 dvss.n1103 dvss.n623 36.1417
R5459 dvss.n1051 dvss.n623 36.1417
R5460 dvss.n1051 dvss.n630 36.1417
R5461 dvss.n1096 dvss.n630 36.1417
R5462 dvss.n1096 dvss.n1095 36.1417
R5463 dvss.n1095 dvss.n1094 36.1417
R5464 dvss.n1094 dvss.n634 36.1417
R5465 dvss.n1088 dvss.n634 36.1417
R5466 dvss.n1088 dvss.n1087 36.1417
R5467 dvss.n1087 dvss.n1086 36.1417
R5468 dvss.n1086 dvss.n643 36.1417
R5469 dvss.n670 dvss.n643 36.1417
R5470 dvss.n670 dvss.n653 36.1417
R5471 dvss.n660 dvss.n653 36.1417
R5472 dvss.n661 dvss.n660 36.1417
R5473 dvss.n669 dvss.n661 36.1417
R5474 dvss.n669 dvss.n665 36.1417
R5475 dvss.n665 dvss.n568 36.1417
R5476 dvss.n1295 dvss.n568 36.1417
R5477 dvss.n1295 dvss.n562 36.1417
R5478 dvss.n1320 dvss.n562 36.1417
R5479 dvss.n1320 dvss.n1319 36.1417
R5480 dvss.n1319 dvss.n564 36.1417
R5481 dvss.n1313 dvss.n564 36.1417
R5482 dvss.n1313 dvss.n553 36.1417
R5483 dvss.n553 dvss.n551 36.1417
R5484 dvss.n1335 dvss.n551 36.1417
R5485 dvss.n1335 dvss.n547 36.1417
R5486 dvss.n1348 dvss.n547 36.1417
R5487 dvss.n1348 dvss.n539 36.1417
R5488 dvss.n1363 dvss.n539 36.1417
R5489 dvss.n1364 dvss.n1363 36.1417
R5490 dvss.n1364 dvss.n536 36.1417
R5491 dvss.n536 dvss.n530 36.1417
R5492 dvss.n1384 dvss.n530 36.1417
R5493 dvss.n1385 dvss.n1384 36.1417
R5494 dvss.n1385 dvss.n526 36.1417
R5495 dvss.n526 dvss.n518 36.1417
R5496 dvss.n523 dvss.n518 36.1417
R5497 dvss.n1405 dvss.n523 36.1417
R5498 dvss.n1405 dvss.n509 36.1417
R5499 dvss.n1578 dvss.n509 36.1417
R5500 dvss.n1578 dvss.n510 36.1417
R5501 dvss.n1420 dvss.n510 36.1417
R5502 dvss.n1421 dvss.n1420 36.1417
R5503 dvss.n1425 dvss.n1421 36.1417
R5504 dvss.n1426 dvss.n1425 36.1417
R5505 dvss.n1491 dvss.n1426 36.1417
R5506 dvss.n1491 dvss.n1430 36.1417
R5507 dvss.n1435 dvss.n1430 36.1417
R5508 dvss.n1498 dvss.n1435 36.1417
R5509 dvss.n1501 dvss.n1498 36.1417
R5510 dvss.n1501 dvss.n1441 36.1417
R5511 dvss.n1446 dvss.n1441 36.1417
R5512 dvss.n1447 dvss.n1446 36.1417
R5513 dvss.n1468 dvss.n1447 36.1417
R5514 dvss.n1468 dvss.n1450 36.1417
R5515 dvss.n1458 dvss.n1450 36.1417
R5516 dvss.n1459 dvss.n1458 36.1417
R5517 dvss.n1467 dvss.n1459 36.1417
R5518 dvss.n1467 dvss.n1463 36.1417
R5519 dvss.n1463 dvss.n458 36.1417
R5520 dvss.n2885 dvss.n458 36.1417
R5521 dvss.n2885 dvss.n453 36.1417
R5522 dvss.n2912 dvss.n453 36.1417
R5523 dvss.n2912 dvss.n454 36.1417
R5524 dvss.n2899 dvss.n454 36.1417
R5525 dvss.n2905 dvss.n2899 36.1417
R5526 dvss.n2905 dvss.n444 36.1417
R5527 dvss.n444 dvss.n442 36.1417
R5528 dvss.n2927 dvss.n442 36.1417
R5529 dvss.n2927 dvss.n438 36.1417
R5530 dvss.n2940 dvss.n438 36.1417
R5531 dvss.n2940 dvss.n430 36.1417
R5532 dvss.n2955 dvss.n430 36.1417
R5533 dvss.n2956 dvss.n2955 36.1417
R5534 dvss.n2956 dvss.n427 36.1417
R5535 dvss.n427 dvss.n421 36.1417
R5536 dvss.n2976 dvss.n421 36.1417
R5537 dvss.n2977 dvss.n2976 36.1417
R5538 dvss.n2977 dvss.n417 36.1417
R5539 dvss.n417 dvss.n409 36.1417
R5540 dvss.n414 dvss.n409 36.1417
R5541 dvss.n2998 dvss.n414 36.1417
R5542 dvss.n2998 dvss.n400 36.1417
R5543 dvss.n3013 dvss.n400 36.1417
R5544 dvss.n3013 dvss.n394 36.1417
R5545 dvss.n3032 dvss.n394 36.1417
R5546 dvss.n3032 dvss.n395 36.1417
R5547 dvss.n395 dvss.n388 36.1417
R5548 dvss.n3038 dvss.n388 36.1417
R5549 dvss.n3038 dvss.n383 36.1417
R5550 dvss.n3049 dvss.n383 36.1417
R5551 dvss.n3049 dvss.n378 36.1417
R5552 dvss.n3058 dvss.n378 36.1417
R5553 dvss.n3058 dvss.n373 36.1417
R5554 dvss.n3075 dvss.n373 36.1417
R5555 dvss.n3075 dvss.n366 36.1417
R5556 dvss.n3082 dvss.n366 36.1417
R5557 dvss.n3082 dvss.n362 36.1417
R5558 dvss.n3092 dvss.n362 36.1417
R5559 dvss.n3092 dvss.n357 36.1417
R5560 dvss.n3106 dvss.n357 36.1417
R5561 dvss.n3106 dvss.n346 36.1417
R5562 dvss.n3115 dvss.n346 36.1417
R5563 dvss.n3115 dvss.n340 36.1417
R5564 dvss.n3127 dvss.n340 36.1417
R5565 dvss.n3128 dvss.n3127 36.1417
R5566 dvss.n3128 dvss.n335 36.1417
R5567 dvss.n335 dvss.n328 36.1417
R5568 dvss.n329 dvss.n328 36.1417
R5569 dvss.n3141 dvss.n329 36.1417
R5570 dvss.n3141 dvss.n320 36.1417
R5571 dvss.n320 dvss.n318 36.1417
R5572 dvss.n3166 dvss.n318 36.1417
R5573 dvss.n3166 dvss.n313 36.1417
R5574 dvss.n3175 dvss.n313 36.1417
R5575 dvss.n3175 dvss.n308 36.1417
R5576 dvss.n3188 dvss.n308 36.1417
R5577 dvss.n3188 dvss.n302 36.1417
R5578 dvss.n3198 dvss.n302 36.1417
R5579 dvss.n3198 dvss.n298 36.1417
R5580 dvss.n3208 dvss.n298 36.1417
R5581 dvss.n3208 dvss.n293 36.1417
R5582 dvss.n3222 dvss.n293 36.1417
R5583 dvss.n3222 dvss.n282 36.1417
R5584 dvss.n3231 dvss.n282 36.1417
R5585 dvss.n3231 dvss.n276 36.1417
R5586 dvss.n3243 dvss.n276 36.1417
R5587 dvss.n3244 dvss.n3243 36.1417
R5588 dvss.n3244 dvss.n271 36.1417
R5589 dvss.n271 dvss.n264 36.1417
R5590 dvss.n265 dvss.n264 36.1417
R5591 dvss.n3257 dvss.n265 36.1417
R5592 dvss.n3257 dvss.n255 36.1417
R5593 dvss.n3275 dvss.n255 36.1417
R5594 dvss.n3276 dvss.n3275 36.1417
R5595 dvss.n3276 dvss.n252 36.1417
R5596 dvss.n252 dvss.n246 36.1417
R5597 dvss.n246 dvss.n241 36.1417
R5598 dvss.n3307 dvss.n241 36.1417
R5599 dvss.n3307 dvss.n242 36.1417
R5600 dvss.n242 dvss.n237 36.1417
R5601 dvss.n237 dvss.n231 36.1417
R5602 dvss.n3324 dvss.n231 36.1417
R5603 dvss.n3325 dvss.n3324 36.1417
R5604 dvss.n3325 dvss.n227 36.1417
R5605 dvss.n227 dvss.n219 36.1417
R5606 dvss.n224 dvss.n219 36.1417
R5607 dvss.n3345 dvss.n224 36.1417
R5608 dvss.n3345 dvss.n210 36.1417
R5609 dvss.n3544 dvss.n210 36.1417
R5610 dvss.n3544 dvss.n211 36.1417
R5611 dvss.n3360 dvss.n211 36.1417
R5612 dvss.n3361 dvss.n3360 36.1417
R5613 dvss.n3365 dvss.n3361 36.1417
R5614 dvss.n3366 dvss.n3365 36.1417
R5615 dvss.n3429 dvss.n3366 36.1417
R5616 dvss.n3429 dvss.n3370 36.1417
R5617 dvss.n3375 dvss.n3370 36.1417
R5618 dvss.n3425 dvss.n3375 36.1417
R5619 dvss.n3428 dvss.n3425 36.1417
R5620 dvss.n3428 dvss.n3381 36.1417
R5621 dvss.n3386 dvss.n3381 36.1417
R5622 dvss.n3387 dvss.n3386 36.1417
R5623 dvss.n3422 dvss.n3387 36.1417
R5624 dvss.n3422 dvss.n3390 36.1417
R5625 dvss.n3395 dvss.n3390 36.1417
R5626 dvss.n3396 dvss.n3395 36.1417
R5627 dvss.n3415 dvss.n3396 36.1417
R5628 dvss.n3476 dvss.n3415 36.1417
R5629 dvss.n3476 dvss.n3416 36.1417
R5630 dvss.n3416 dvss.n3411 36.1417
R5631 dvss.n3411 dvss.n3405 36.1417
R5632 dvss.n3409 dvss.n3405 36.1417
R5633 dvss.n3489 dvss.n3409 36.1417
R5634 dvss.n3489 dvss.n125 36.1417
R5635 dvss.n854 dvss.n853 36.1417
R5636 dvss.n853 dvss.n852 36.1417
R5637 dvss.n852 dvss.n771 36.1417
R5638 dvss.n775 dvss.n771 36.1417
R5639 dvss.n845 dvss.n775 36.1417
R5640 dvss.n845 dvss.n844 36.1417
R5641 dvss.n844 dvss.n843 36.1417
R5642 dvss.n843 dvss.n779 36.1417
R5643 dvss.n837 dvss.n779 36.1417
R5644 dvss.n837 dvss.n836 36.1417
R5645 dvss.n836 dvss.n835 36.1417
R5646 dvss.n835 dvss.n804 36.1417
R5647 dvss.n829 dvss.n804 36.1417
R5648 dvss.n829 dvss.n828 36.1417
R5649 dvss.n828 dvss.n827 36.1417
R5650 dvss.n827 dvss.n821 36.1417
R5651 dvss.n821 dvss.n611 36.1417
R5652 dvss.n1113 dvss.n611 36.1417
R5653 dvss.n1113 dvss.n610 36.1417
R5654 dvss.n1118 dvss.n610 36.1417
R5655 dvss.n1118 dvss.n607 36.1417
R5656 dvss.n1124 dvss.n607 36.1417
R5657 dvss.n1124 dvss.n606 36.1417
R5658 dvss.n1130 dvss.n606 36.1417
R5659 dvss.n1130 dvss.n602 36.1417
R5660 dvss.n1136 dvss.n602 36.1417
R5661 dvss.n1136 dvss.n598 36.1417
R5662 dvss.n1145 dvss.n598 36.1417
R5663 dvss.n1145 dvss.n594 36.1417
R5664 dvss.n1152 dvss.n594 36.1417
R5665 dvss.n1152 dvss.n588 36.1417
R5666 dvss.n1160 dvss.n588 36.1417
R5667 dvss.n1160 dvss.n585 36.1417
R5668 dvss.n1167 dvss.n585 36.1417
R5669 dvss.n1167 dvss.n580 36.1417
R5670 dvss.n1175 dvss.n580 36.1417
R5671 dvss.n1175 dvss.n577 36.1417
R5672 dvss.n1181 dvss.n577 36.1417
R5673 dvss.n1181 dvss.n575 36.1417
R5674 dvss.n1288 dvss.n575 36.1417
R5675 dvss.n1288 dvss.n576 36.1417
R5676 dvss.n1284 dvss.n576 36.1417
R5677 dvss.n1284 dvss.n1283 36.1417
R5678 dvss.n1283 dvss.n1186 36.1417
R5679 dvss.n1279 dvss.n1186 36.1417
R5680 dvss.n1279 dvss.n1278 36.1417
R5681 dvss.n1278 dvss.n1189 36.1417
R5682 dvss.n1192 dvss.n1189 36.1417
R5683 dvss.n1270 dvss.n1192 36.1417
R5684 dvss.n1270 dvss.n1269 36.1417
R5685 dvss.n1269 dvss.n1195 36.1417
R5686 dvss.n1261 dvss.n1195 36.1417
R5687 dvss.n1261 dvss.n1260 36.1417
R5688 dvss.n1260 dvss.n1201 36.1417
R5689 dvss.n1253 dvss.n1201 36.1417
R5690 dvss.n1253 dvss.n1252 36.1417
R5691 dvss.n1252 dvss.n1205 36.1417
R5692 dvss.n1209 dvss.n1205 36.1417
R5693 dvss.n1243 dvss.n1209 36.1417
R5694 dvss.n1243 dvss.n1242 36.1417
R5695 dvss.n1242 dvss.n501 36.1417
R5696 dvss.n1586 dvss.n501 36.1417
R5697 dvss.n1586 dvss.n500 36.1417
R5698 dvss.n1591 dvss.n500 36.1417
R5699 dvss.n1591 dvss.n497 36.1417
R5700 dvss.n1597 dvss.n497 36.1417
R5701 dvss.n1597 dvss.n496 36.1417
R5702 dvss.n1603 dvss.n496 36.1417
R5703 dvss.n1603 dvss.n492 36.1417
R5704 dvss.n1609 dvss.n492 36.1417
R5705 dvss.n1609 dvss.n488 36.1417
R5706 dvss.n1618 dvss.n488 36.1417
R5707 dvss.n1618 dvss.n484 36.1417
R5708 dvss.n1625 dvss.n484 36.1417
R5709 dvss.n1625 dvss.n478 36.1417
R5710 dvss.n1633 dvss.n478 36.1417
R5711 dvss.n1633 dvss.n475 36.1417
R5712 dvss.n1640 dvss.n475 36.1417
R5713 dvss.n1640 dvss.n470 36.1417
R5714 dvss.n1648 dvss.n470 36.1417
R5715 dvss.n1648 dvss.n467 36.1417
R5716 dvss.n1654 dvss.n467 36.1417
R5717 dvss.n1654 dvss.n465 36.1417
R5718 dvss.n2878 dvss.n465 36.1417
R5719 dvss.n2878 dvss.n466 36.1417
R5720 dvss.n2874 dvss.n466 36.1417
R5721 dvss.n2874 dvss.n2873 36.1417
R5722 dvss.n2873 dvss.n1659 36.1417
R5723 dvss.n2869 dvss.n1659 36.1417
R5724 dvss.n2869 dvss.n2868 36.1417
R5725 dvss.n2868 dvss.n1662 36.1417
R5726 dvss.n1665 dvss.n1662 36.1417
R5727 dvss.n2860 dvss.n1665 36.1417
R5728 dvss.n2860 dvss.n2859 36.1417
R5729 dvss.n2859 dvss.n1668 36.1417
R5730 dvss.n2851 dvss.n1668 36.1417
R5731 dvss.n2851 dvss.n2850 36.1417
R5732 dvss.n2850 dvss.n1674 36.1417
R5733 dvss.n2843 dvss.n1674 36.1417
R5734 dvss.n2843 dvss.n2842 36.1417
R5735 dvss.n2842 dvss.n1678 36.1417
R5736 dvss.n1682 dvss.n1678 36.1417
R5737 dvss.n2833 dvss.n1682 36.1417
R5738 dvss.n2833 dvss.n2832 36.1417
R5739 dvss.n2832 dvss.n1685 36.1417
R5740 dvss.n2828 dvss.n1685 36.1417
R5741 dvss.n2828 dvss.n2827 36.1417
R5742 dvss.n2827 dvss.n1688 36.1417
R5743 dvss.n2823 dvss.n1688 36.1417
R5744 dvss.n2823 dvss.n2822 36.1417
R5745 dvss.n2822 dvss.n1691 36.1417
R5746 dvss.n2818 dvss.n1691 36.1417
R5747 dvss.n2818 dvss.n2817 36.1417
R5748 dvss.n2817 dvss.n1694 36.1417
R5749 dvss.n2810 dvss.n1694 36.1417
R5750 dvss.n2810 dvss.n2809 36.1417
R5751 dvss.n2809 dvss.n1699 36.1417
R5752 dvss.n2801 dvss.n1699 36.1417
R5753 dvss.n2801 dvss.n2800 36.1417
R5754 dvss.n2800 dvss.n1705 36.1417
R5755 dvss.n2793 dvss.n1705 36.1417
R5756 dvss.n2793 dvss.n2792 36.1417
R5757 dvss.n2792 dvss.n1709 36.1417
R5758 dvss.n1713 dvss.n1709 36.1417
R5759 dvss.n2783 dvss.n1713 36.1417
R5760 dvss.n2783 dvss.n2782 36.1417
R5761 dvss.n2782 dvss.n1716 36.1417
R5762 dvss.n2778 dvss.n1716 36.1417
R5763 dvss.n2778 dvss.n2777 36.1417
R5764 dvss.n2777 dvss.n1719 36.1417
R5765 dvss.n2773 dvss.n1719 36.1417
R5766 dvss.n2773 dvss.n2772 36.1417
R5767 dvss.n2772 dvss.n1722 36.1417
R5768 dvss.n2768 dvss.n1722 36.1417
R5769 dvss.n2768 dvss.n2767 36.1417
R5770 dvss.n2767 dvss.n1725 36.1417
R5771 dvss.n2760 dvss.n1725 36.1417
R5772 dvss.n2760 dvss.n2759 36.1417
R5773 dvss.n2759 dvss.n1730 36.1417
R5774 dvss.n2751 dvss.n1730 36.1417
R5775 dvss.n2751 dvss.n2750 36.1417
R5776 dvss.n2750 dvss.n1736 36.1417
R5777 dvss.n2743 dvss.n1736 36.1417
R5778 dvss.n2743 dvss.n2742 36.1417
R5779 dvss.n2742 dvss.n1740 36.1417
R5780 dvss.n1744 dvss.n1740 36.1417
R5781 dvss.n2733 dvss.n1744 36.1417
R5782 dvss.n2733 dvss.n2732 36.1417
R5783 dvss.n2732 dvss.n1747 36.1417
R5784 dvss.n2728 dvss.n1747 36.1417
R5785 dvss.n2728 dvss.n2727 36.1417
R5786 dvss.n2727 dvss.n1750 36.1417
R5787 dvss.n2723 dvss.n1750 36.1417
R5788 dvss.n2723 dvss.n2722 36.1417
R5789 dvss.n2722 dvss.n1753 36.1417
R5790 dvss.n2718 dvss.n1753 36.1417
R5791 dvss.n2718 dvss.n2717 36.1417
R5792 dvss.n2717 dvss.n1756 36.1417
R5793 dvss.n2710 dvss.n1756 36.1417
R5794 dvss.n2710 dvss.n2709 36.1417
R5795 dvss.n2709 dvss.n1761 36.1417
R5796 dvss.n2701 dvss.n1761 36.1417
R5797 dvss.n2701 dvss.n2700 36.1417
R5798 dvss.n2700 dvss.n1767 36.1417
R5799 dvss.n2693 dvss.n1767 36.1417
R5800 dvss.n2693 dvss.n2692 36.1417
R5801 dvss.n2692 dvss.n1771 36.1417
R5802 dvss.n1776 dvss.n1771 36.1417
R5803 dvss.n2683 dvss.n1776 36.1417
R5804 dvss.n2683 dvss.n168 36.1417
R5805 dvss.n3551 dvss.n168 36.1417
R5806 dvss.n3551 dvss.n166 36.1417
R5807 dvss.n3568 dvss.n166 36.1417
R5808 dvss.n3568 dvss.n167 36.1417
R5809 dvss.n3564 dvss.n167 36.1417
R5810 dvss.n3564 dvss.n3563 36.1417
R5811 dvss.n3563 dvss.n3559 36.1417
R5812 dvss.n3559 dvss.n160 36.1417
R5813 dvss.n3576 dvss.n160 36.1417
R5814 dvss.n3576 dvss.n157 36.1417
R5815 dvss.n3587 dvss.n157 36.1417
R5816 dvss.n3587 dvss.n154 36.1417
R5817 dvss.n3593 dvss.n154 36.1417
R5818 dvss.n3593 dvss.n149 36.1417
R5819 dvss.n3602 dvss.n149 36.1417
R5820 dvss.n3602 dvss.n144 36.1417
R5821 dvss.n3608 dvss.n144 36.1417
R5822 dvss.n3608 dvss.n143 36.1417
R5823 dvss.n3620 dvss.n143 36.1417
R5824 dvss.n3620 dvss.n139 36.1417
R5825 dvss.n3626 dvss.n139 36.1417
R5826 dvss.n3626 dvss.n137 36.1417
R5827 dvss.n3633 dvss.n137 36.1417
R5828 dvss.n3633 dvss.n138 36.1417
R5829 dvss.n138 dvss.n133 36.1417
R5830 dvss.n133 dvss.n131 36.1417
R5831 dvss.n3642 dvss.n131 36.1417
R5832 dvss.n956 dvss.n861 36.1417
R5833 dvss.n957 dvss.n956 36.1417
R5834 dvss.n957 dvss.n761 36.1417
R5835 dvss.n966 dvss.n761 36.1417
R5836 dvss.n966 dvss.n753 36.1417
R5837 dvss.n979 dvss.n753 36.1417
R5838 dvss.n979 dvss.n746 36.1417
R5839 dvss.n992 dvss.n746 36.1417
R5840 dvss.n992 dvss.n741 36.1417
R5841 dvss.n1001 dvss.n741 36.1417
R5842 dvss.n1001 dvss.n735 36.1417
R5843 dvss.n1017 dvss.n735 36.1417
R5844 dvss.n1017 dvss.n726 36.1417
R5845 dvss.n1032 dvss.n726 36.1417
R5846 dvss.n1032 dvss.n1031 36.1417
R5847 dvss.n1031 dvss.n718 36.1417
R5848 dvss.n1041 dvss.n718 36.1417
R5849 dvss.n1042 dvss.n1041 36.1417
R5850 dvss.n1043 dvss.n1042 36.1417
R5851 dvss.n1043 dvss.n714 36.1417
R5852 dvss.n1048 dvss.n714 36.1417
R5853 dvss.n1059 dvss.n712 36.1417
R5854 dvss.n1060 dvss.n1059 36.1417
R5855 dvss.n1063 dvss.n1060 36.1417
R5856 dvss.n1064 dvss.n1063 36.1417
R5857 dvss.n1066 dvss.n1064 36.1417
R5858 dvss.n1066 dvss.n1065 36.1417
R5859 dvss.n1065 dvss.n649 36.1417
R5860 dvss.n1082 dvss.n649 36.1417
R5861 dvss.n1082 dvss.n1081 36.1417
R5862 dvss.n1081 dvss.n650 36.1417
R5863 dvss.n706 dvss.n650 36.1417
R5864 dvss.n706 dvss.n705 36.1417
R5865 dvss.n705 dvss.n656 36.1417
R5866 dvss.n666 dvss.n656 36.1417
R5867 dvss.n692 dvss.n666 36.1417
R5868 dvss.n692 dvss.n691 36.1417
R5869 dvss.n691 dvss.n565 36.1417
R5870 dvss.n1301 dvss.n565 36.1417
R5871 dvss.n1302 dvss.n1301 36.1417
R5872 dvss.n1317 dvss.n1302 36.1417
R5873 dvss.n1317 dvss.n1316 36.1417
R5874 dvss.n1327 dvss.n554 36.1417
R5875 dvss.n1327 dvss.n1326 36.1417
R5876 dvss.n1326 dvss.n548 36.1417
R5877 dvss.n1340 dvss.n548 36.1417
R5878 dvss.n1340 dvss.n542 36.1417
R5879 dvss.n1353 dvss.n542 36.1417
R5880 dvss.n1353 dvss.n538 36.1417
R5881 dvss.n1367 dvss.n538 36.1417
R5882 dvss.n1367 dvss.n533 36.1417
R5883 dvss.n1377 dvss.n533 36.1417
R5884 dvss.n1377 dvss.n529 36.1417
R5885 dvss.n1394 dvss.n529 36.1417
R5886 dvss.n1394 dvss.n520 36.1417
R5887 dvss.n1409 dvss.n520 36.1417
R5888 dvss.n1409 dvss.n1408 36.1417
R5889 dvss.n1408 dvss.n512 36.1417
R5890 dvss.n1417 dvss.n512 36.1417
R5891 dvss.n1576 dvss.n1417 36.1417
R5892 dvss.n1576 dvss.n1575 36.1417
R5893 dvss.n1575 dvss.n1419 36.1417
R5894 dvss.n1571 dvss.n1419 36.1417
R5895 dvss.n1570 dvss.n1424 36.1417
R5896 dvss.n1431 dvss.n1424 36.1417
R5897 dvss.n1563 dvss.n1431 36.1417
R5898 dvss.n1563 dvss.n1562 36.1417
R5899 dvss.n1562 dvss.n1434 36.1417
R5900 dvss.n1442 dvss.n1434 36.1417
R5901 dvss.n1554 dvss.n1442 36.1417
R5902 dvss.n1554 dvss.n1553 36.1417
R5903 dvss.n1553 dvss.n1445 36.1417
R5904 dvss.n1451 dvss.n1445 36.1417
R5905 dvss.n1543 dvss.n1451 36.1417
R5906 dvss.n1543 dvss.n1542 36.1417
R5907 dvss.n1542 dvss.n1454 36.1417
R5908 dvss.n1464 dvss.n1454 36.1417
R5909 dvss.n1529 dvss.n1464 36.1417
R5910 dvss.n1529 dvss.n1528 36.1417
R5911 dvss.n1528 dvss.n455 36.1417
R5912 dvss.n2891 dvss.n455 36.1417
R5913 dvss.n2910 dvss.n2891 36.1417
R5914 dvss.n2910 dvss.n2909 36.1417
R5915 dvss.n2909 dvss.n2898 36.1417
R5916 dvss.n2919 dvss.n445 36.1417
R5917 dvss.n2919 dvss.n2918 36.1417
R5918 dvss.n2918 dvss.n439 36.1417
R5919 dvss.n2932 dvss.n439 36.1417
R5920 dvss.n2932 dvss.n433 36.1417
R5921 dvss.n2945 dvss.n433 36.1417
R5922 dvss.n2945 dvss.n429 36.1417
R5923 dvss.n2959 dvss.n429 36.1417
R5924 dvss.n2959 dvss.n424 36.1417
R5925 dvss.n2969 dvss.n424 36.1417
R5926 dvss.n2969 dvss.n420 36.1417
R5927 dvss.n2986 dvss.n420 36.1417
R5928 dvss.n2986 dvss.n411 36.1417
R5929 dvss.n3002 dvss.n411 36.1417
R5930 dvss.n3002 dvss.n3001 36.1417
R5931 dvss.n3001 dvss.n403 36.1417
R5932 dvss.n3010 dvss.n403 36.1417
R5933 dvss.n3011 dvss.n3010 36.1417
R5934 dvss.n3011 dvss.n396 36.1417
R5935 dvss.n3030 dvss.n396 36.1417
R5936 dvss.n3030 dvss.n3029 36.1417
R5937 dvss.n3026 dvss.n386 36.1417
R5938 dvss.n3046 dvss.n386 36.1417
R5939 dvss.n3047 dvss.n3046 36.1417
R5940 dvss.n3047 dvss.n381 36.1417
R5941 dvss.n381 dvss.n374 36.1417
R5942 dvss.n3072 dvss.n374 36.1417
R5943 dvss.n3073 dvss.n3072 36.1417
R5944 dvss.n3073 dvss.n364 36.1417
R5945 dvss.n3084 dvss.n364 36.1417
R5946 dvss.n3085 dvss.n3084 36.1417
R5947 dvss.n3085 dvss.n358 36.1417
R5948 dvss.n3097 dvss.n358 36.1417
R5949 dvss.n3097 dvss.n348 36.1417
R5950 dvss.n3119 dvss.n348 36.1417
R5951 dvss.n3119 dvss.n3118 36.1417
R5952 dvss.n3118 dvss.n351 36.1417
R5953 dvss.n351 dvss.n338 36.1417
R5954 dvss.n3131 dvss.n338 36.1417
R5955 dvss.n3131 dvss.n326 36.1417
R5956 dvss.n3145 dvss.n326 36.1417
R5957 dvss.n3145 dvss.n327 36.1417
R5958 dvss.n3152 dvss.n321 36.1417
R5959 dvss.n3152 dvss.n3151 36.1417
R5960 dvss.n3151 dvss.n316 36.1417
R5961 dvss.n316 dvss.n311 36.1417
R5962 dvss.n3177 dvss.n311 36.1417
R5963 dvss.n3178 dvss.n3177 36.1417
R5964 dvss.n3178 dvss.n306 36.1417
R5965 dvss.n306 dvss.n300 36.1417
R5966 dvss.n3200 dvss.n300 36.1417
R5967 dvss.n3201 dvss.n3200 36.1417
R5968 dvss.n3201 dvss.n294 36.1417
R5969 dvss.n3213 dvss.n294 36.1417
R5970 dvss.n3213 dvss.n284 36.1417
R5971 dvss.n3235 dvss.n284 36.1417
R5972 dvss.n3235 dvss.n3234 36.1417
R5973 dvss.n3234 dvss.n287 36.1417
R5974 dvss.n287 dvss.n274 36.1417
R5975 dvss.n3247 dvss.n274 36.1417
R5976 dvss.n3247 dvss.n262 36.1417
R5977 dvss.n3261 dvss.n262 36.1417
R5978 dvss.n3261 dvss.n263 36.1417
R5979 dvss.n3267 dvss.n257 36.1417
R5980 dvss.n3267 dvss.n254 36.1417
R5981 dvss.n3284 dvss.n254 36.1417
R5982 dvss.n3284 dvss.n247 36.1417
R5983 dvss.n3292 dvss.n247 36.1417
R5984 dvss.n3292 dvss.n243 36.1417
R5985 dvss.n3305 dvss.n243 36.1417
R5986 dvss.n3305 dvss.n3304 36.1417
R5987 dvss.n3304 dvss.n234 36.1417
R5988 dvss.n3317 dvss.n234 36.1417
R5989 dvss.n3317 dvss.n230 36.1417
R5990 dvss.n3334 dvss.n230 36.1417
R5991 dvss.n3334 dvss.n221 36.1417
R5992 dvss.n3349 dvss.n221 36.1417
R5993 dvss.n3349 dvss.n3348 36.1417
R5994 dvss.n3348 dvss.n213 36.1417
R5995 dvss.n3357 dvss.n213 36.1417
R5996 dvss.n3542 dvss.n3357 36.1417
R5997 dvss.n3542 dvss.n3541 36.1417
R5998 dvss.n3541 dvss.n3359 36.1417
R5999 dvss.n3537 dvss.n3359 36.1417
R6000 dvss.n3536 dvss.n3364 36.1417
R6001 dvss.n3371 dvss.n3364 36.1417
R6002 dvss.n3529 dvss.n3371 36.1417
R6003 dvss.n3529 dvss.n3528 36.1417
R6004 dvss.n3528 dvss.n3374 36.1417
R6005 dvss.n3382 dvss.n3374 36.1417
R6006 dvss.n3520 dvss.n3382 36.1417
R6007 dvss.n3520 dvss.n3519 36.1417
R6008 dvss.n3519 dvss.n3385 36.1417
R6009 dvss.n3391 dvss.n3385 36.1417
R6010 dvss.n3509 dvss.n3391 36.1417
R6011 dvss.n3509 dvss.n3508 36.1417
R6012 dvss.n3508 dvss.n3394 36.1417
R6013 dvss.n3473 dvss.n3394 36.1417
R6014 dvss.n3474 dvss.n3473 36.1417
R6015 dvss.n3474 dvss.n3413 36.1417
R6016 dvss.n3413 dvss.n3406 36.1417
R6017 dvss.n3493 dvss.n3406 36.1417
R6018 dvss.n3493 dvss.n3492 36.1417
R6019 dvss.n3492 dvss.n124 36.1417
R6020 dvss.n3647 dvss.n124 36.1417
R6021 dvss.n2664 dvss.n1966 36.1417
R6022 dvss.n2661 dvss.n1966 36.1417
R6023 dvss.n2661 dvss.n2660 36.1417
R6024 dvss.n2660 dvss.n1969 36.1417
R6025 dvss.n2655 dvss.n1969 36.1417
R6026 dvss.n2655 dvss.n2654 36.1417
R6027 dvss.n2654 dvss.n1974 36.1417
R6028 dvss.n2650 dvss.n1974 36.1417
R6029 dvss.n2650 dvss.n2649 36.1417
R6030 dvss.n2649 dvss.n1977 36.1417
R6031 dvss.n2642 dvss.n1977 36.1417
R6032 dvss.n2642 dvss.n2641 36.1417
R6033 dvss.n2641 dvss.n1985 36.1417
R6034 dvss.n1990 dvss.n1985 36.1417
R6035 dvss.n2634 dvss.n1990 36.1417
R6036 dvss.n2634 dvss.n2633 36.1417
R6037 dvss.n2630 dvss.n2629 36.1417
R6038 dvss.n2629 dvss.n1997 36.1417
R6039 dvss.n2623 dvss.n1997 36.1417
R6040 dvss.n2623 dvss.n2622 36.1417
R6041 dvss.n2622 dvss.n2003 36.1417
R6042 dvss.n2618 dvss.n2003 36.1417
R6043 dvss.n2618 dvss.n2617 36.1417
R6044 dvss.n2617 dvss.n2008 36.1417
R6045 dvss.n2613 dvss.n2008 36.1417
R6046 dvss.n2613 dvss.n2612 36.1417
R6047 dvss.n2612 dvss.n2011 36.1417
R6048 dvss.n2605 dvss.n2011 36.1417
R6049 dvss.n2605 dvss.n2604 36.1417
R6050 dvss.n2604 dvss.n2018 36.1417
R6051 dvss.n2597 dvss.n2018 36.1417
R6052 dvss.n2597 dvss.n2596 36.1417
R6053 dvss.n2596 dvss.n2022 36.1417
R6054 dvss.n2589 dvss.n2022 36.1417
R6055 dvss.n2589 dvss.n2588 36.1417
R6056 dvss.n2588 dvss.n2027 36.1417
R6057 dvss.n2584 dvss.n2027 36.1417
R6058 dvss.n2583 dvss.n2030 36.1417
R6059 dvss.n2036 dvss.n2030 36.1417
R6060 dvss.n2576 dvss.n2036 36.1417
R6061 dvss.n2576 dvss.n2575 36.1417
R6062 dvss.n2575 dvss.n2039 36.1417
R6063 dvss.n2571 dvss.n2039 36.1417
R6064 dvss.n2571 dvss.n2570 36.1417
R6065 dvss.n2570 dvss.n2044 36.1417
R6066 dvss.n2566 dvss.n2044 36.1417
R6067 dvss.n2566 dvss.n2565 36.1417
R6068 dvss.n2565 dvss.n2047 36.1417
R6069 dvss.n2558 dvss.n2047 36.1417
R6070 dvss.n2558 dvss.n2557 36.1417
R6071 dvss.n2557 dvss.n2054 36.1417
R6072 dvss.n2550 dvss.n2054 36.1417
R6073 dvss.n2550 dvss.n2549 36.1417
R6074 dvss.n2549 dvss.n2058 36.1417
R6075 dvss.n2542 dvss.n2058 36.1417
R6076 dvss.n2542 dvss.n2541 36.1417
R6077 dvss.n2541 dvss.n2063 36.1417
R6078 dvss.n2537 dvss.n2063 36.1417
R6079 dvss.n2536 dvss.n2066 36.1417
R6080 dvss.n2072 dvss.n2066 36.1417
R6081 dvss.n2529 dvss.n2072 36.1417
R6082 dvss.n2529 dvss.n2528 36.1417
R6083 dvss.n2528 dvss.n2075 36.1417
R6084 dvss.n2524 dvss.n2075 36.1417
R6085 dvss.n2524 dvss.n2523 36.1417
R6086 dvss.n2523 dvss.n2080 36.1417
R6087 dvss.n2519 dvss.n2080 36.1417
R6088 dvss.n2519 dvss.n2518 36.1417
R6089 dvss.n2518 dvss.n2083 36.1417
R6090 dvss.n2511 dvss.n2083 36.1417
R6091 dvss.n2511 dvss.n2510 36.1417
R6092 dvss.n2510 dvss.n2090 36.1417
R6093 dvss.n2503 dvss.n2090 36.1417
R6094 dvss.n2503 dvss.n2502 36.1417
R6095 dvss.n2502 dvss.n2094 36.1417
R6096 dvss.n2495 dvss.n2094 36.1417
R6097 dvss.n2495 dvss.n2494 36.1417
R6098 dvss.n2494 dvss.n2099 36.1417
R6099 dvss.n2490 dvss.n2099 36.1417
R6100 dvss.n2489 dvss.n2102 36.1417
R6101 dvss.n2108 dvss.n2102 36.1417
R6102 dvss.n2482 dvss.n2108 36.1417
R6103 dvss.n2482 dvss.n2481 36.1417
R6104 dvss.n2481 dvss.n2111 36.1417
R6105 dvss.n2477 dvss.n2111 36.1417
R6106 dvss.n2477 dvss.n2476 36.1417
R6107 dvss.n2476 dvss.n2116 36.1417
R6108 dvss.n2472 dvss.n2116 36.1417
R6109 dvss.n2472 dvss.n2471 36.1417
R6110 dvss.n2471 dvss.n2119 36.1417
R6111 dvss.n2464 dvss.n2119 36.1417
R6112 dvss.n2464 dvss.n2463 36.1417
R6113 dvss.n2463 dvss.n2126 36.1417
R6114 dvss.n2456 dvss.n2126 36.1417
R6115 dvss.n2456 dvss.n2455 36.1417
R6116 dvss.n2455 dvss.n2130 36.1417
R6117 dvss.n2448 dvss.n2130 36.1417
R6118 dvss.n2448 dvss.n2447 36.1417
R6119 dvss.n2447 dvss.n2135 36.1417
R6120 dvss.n2443 dvss.n2135 36.1417
R6121 dvss.n2442 dvss.n2138 36.1417
R6122 dvss.n2144 dvss.n2138 36.1417
R6123 dvss.n2435 dvss.n2144 36.1417
R6124 dvss.n2435 dvss.n2434 36.1417
R6125 dvss.n2434 dvss.n2147 36.1417
R6126 dvss.n2430 dvss.n2147 36.1417
R6127 dvss.n2430 dvss.n2429 36.1417
R6128 dvss.n2429 dvss.n2152 36.1417
R6129 dvss.n2425 dvss.n2152 36.1417
R6130 dvss.n2425 dvss.n2424 36.1417
R6131 dvss.n2424 dvss.n2155 36.1417
R6132 dvss.n2417 dvss.n2155 36.1417
R6133 dvss.n2417 dvss.n2416 36.1417
R6134 dvss.n2416 dvss.n2162 36.1417
R6135 dvss.n2409 dvss.n2162 36.1417
R6136 dvss.n2409 dvss.n2408 36.1417
R6137 dvss.n2408 dvss.n2166 36.1417
R6138 dvss.n2401 dvss.n2166 36.1417
R6139 dvss.n2401 dvss.n2400 36.1417
R6140 dvss.n2400 dvss.n2171 36.1417
R6141 dvss.n2396 dvss.n2171 36.1417
R6142 dvss.n2395 dvss.n2174 36.1417
R6143 dvss.n2180 dvss.n2174 36.1417
R6144 dvss.n2388 dvss.n2180 36.1417
R6145 dvss.n2388 dvss.n2387 36.1417
R6146 dvss.n2387 dvss.n2183 36.1417
R6147 dvss.n2383 dvss.n2183 36.1417
R6148 dvss.n2383 dvss.n2382 36.1417
R6149 dvss.n2382 dvss.n2188 36.1417
R6150 dvss.n2378 dvss.n2188 36.1417
R6151 dvss.n2378 dvss.n2377 36.1417
R6152 dvss.n2377 dvss.n2192 36.1417
R6153 dvss.n2370 dvss.n2192 36.1417
R6154 dvss.n2370 dvss.n2369 36.1417
R6155 dvss.n2369 dvss.n2196 36.1417
R6156 dvss.n2362 dvss.n2196 36.1417
R6157 dvss.n2362 dvss.n2361 36.1417
R6158 dvss.n2361 dvss.n2200 36.1417
R6159 dvss.n2354 dvss.n2200 36.1417
R6160 dvss.n2354 dvss.n2353 36.1417
R6161 dvss.n2353 dvss.n2203 36.1417
R6162 dvss.n2349 dvss.n2203 36.1417
R6163 dvss.n2348 dvss.n2206 36.1417
R6164 dvss.n2210 dvss.n2206 36.1417
R6165 dvss.n2341 dvss.n2210 36.1417
R6166 dvss.n2341 dvss.n2340 36.1417
R6167 dvss.n2340 dvss.n2213 36.1417
R6168 dvss.n2336 dvss.n2213 36.1417
R6169 dvss.n2336 dvss.n2335 36.1417
R6170 dvss.n2335 dvss.n2216 36.1417
R6171 dvss.n2331 dvss.n2216 36.1417
R6172 dvss.n2331 dvss.n2330 36.1417
R6173 dvss.n2330 dvss.n2246 36.1417
R6174 dvss.n2323 dvss.n2246 36.1417
R6175 dvss.n2323 dvss.n2322 36.1417
R6176 dvss.n2322 dvss.n2251 36.1417
R6177 dvss.n2315 dvss.n2251 36.1417
R6178 dvss.n2315 dvss.n2314 36.1417
R6179 dvss.n2314 dvss.n2255 36.1417
R6180 dvss.n2307 dvss.n2255 36.1417
R6181 dvss.n2307 dvss.n2306 36.1417
R6182 dvss.n2306 dvss.n2258 36.1417
R6183 dvss.n2302 dvss.n2258 36.1417
R6184 dvss.n2301 dvss.n2292 36.1417
R6185 dvss.n2292 dvss.n68 36.1417
R6186 dvss.n3739 dvss.n68 36.1417
R6187 dvss.n3739 dvss.n3738 36.1417
R6188 dvss.n3738 dvss.n71 36.1417
R6189 dvss.n3734 dvss.n71 36.1417
R6190 dvss.n3734 dvss.n3733 36.1417
R6191 dvss.n3733 dvss.n74 36.1417
R6192 dvss.n3729 dvss.n74 36.1417
R6193 dvss.n3729 dvss.n3728 36.1417
R6194 dvss.n3728 dvss.n77 36.1417
R6195 dvss.n3721 dvss.n77 36.1417
R6196 dvss.n3721 dvss.n3720 36.1417
R6197 dvss.n3720 dvss.n82 36.1417
R6198 dvss.n3713 dvss.n82 36.1417
R6199 dvss.n3713 dvss.n3712 36.1417
R6200 dvss.n3712 dvss.n86 36.1417
R6201 dvss.n3705 dvss.n86 36.1417
R6202 dvss.n3705 dvss.n3704 36.1417
R6203 dvss.n3704 dvss.n89 36.1417
R6204 dvss.n3700 dvss.n89 36.1417
R6205 dvss.n3699 dvss.n92 36.1417
R6206 dvss.n96 dvss.n92 36.1417
R6207 dvss.n3692 dvss.n96 36.1417
R6208 dvss.n3692 dvss.n3691 36.1417
R6209 dvss.n3691 dvss.n99 36.1417
R6210 dvss.n3687 dvss.n99 36.1417
R6211 dvss.n3687 dvss.n3686 36.1417
R6212 dvss.n3686 dvss.n102 36.1417
R6213 dvss.n3682 dvss.n102 36.1417
R6214 dvss.n3682 dvss.n3681 36.1417
R6215 dvss.n3681 dvss.n105 36.1417
R6216 dvss.n3674 dvss.n105 36.1417
R6217 dvss.n3674 dvss.n3673 36.1417
R6218 dvss.n3673 dvss.n110 36.1417
R6219 dvss.n3666 dvss.n110 36.1417
R6220 dvss.n3666 dvss.n3665 36.1417
R6221 dvss.n3665 dvss.n114 36.1417
R6222 dvss.n3658 dvss.n114 36.1417
R6223 dvss.n3658 dvss.n3657 36.1417
R6224 dvss.n3657 dvss.n117 36.1417
R6225 dvss.n3653 dvss.n117 36.1417
R6226 dvss.n2667 dvss.n1894 35.9189
R6227 dvss.n2264 dvss.t135 35.9189
R6228 dvss.t300 dvss.n3420 34.5917
R6229 dvss.t501 dvss.n228 34.5917
R6230 dvss.t224 dvss.n290 34.5917
R6231 dvss.t390 dvss.n354 34.5917
R6232 dvss.t189 dvss.n418 34.5917
R6233 dvss.n1517 dvss.t334 34.5917
R6234 dvss.t408 dvss.n527 34.5917
R6235 dvss.n680 dvss.t424 34.5917
R6236 dvss.t328 dvss.n733 34.5917
R6237 dvss.n3504 dvss 33.9483
R6238 dvss.n3330 dvss 33.9483
R6239 dvss.n3219 dvss 33.9483
R6240 dvss.n3103 dvss 33.9483
R6241 dvss.n2982 dvss 33.9483
R6242 dvss.n1538 dvss 33.9483
R6243 dvss.n1390 dvss 33.9483
R6244 dvss.n701 dvss 33.9483
R6245 dvss.n1013 dvss 33.9483
R6246 dvss.n3617 dvss 33.9483
R6247 dvss.n2688 dvss 33.9483
R6248 dvss.n2738 dvss 33.9483
R6249 dvss.n2788 dvss 33.9483
R6250 dvss.n2838 dvss 33.9483
R6251 dvss.n1644 dvss 33.9483
R6252 dvss.n1248 dvss 33.9483
R6253 dvss.n1171 dvss 33.9483
R6254 dvss.n815 dvss 33.9483
R6255 dvss.n1890 dvss.t497 32.1345
R6256 dvss.n177 dvss.t101 32.1345
R6257 dvss.t109 dvss.n196 31.6138
R6258 dvss.t103 dvss.t294 31.1326
R6259 dvss.t509 dvss.t489 31.1326
R6260 dvss.t139 dvss.t232 31.1326
R6261 dvss.t536 dvss.t396 31.1326
R6262 dvss.t187 dvss.t208 31.1326
R6263 dvss.t340 dvss.t263 31.1326
R6264 dvss.t406 dvss.t517 31.1326
R6265 dvss.t422 dvss.t86 31.1326
R6266 dvss.t326 dvss.t76 31.1326
R6267 dvss.n915 dvss.n914 30.6481
R6268 dvss.t487 dvss.n2670 28.7399
R6269 dvss.t99 dvss.n180 28.7399
R6270 dvss.n93 dvss.t457 28.1205
R6271 dvss.n2293 dvss.t387 28.1205
R6272 dvss.n2207 dvss.t433 28.1205
R6273 dvss.n2175 dvss.t450 28.1205
R6274 dvss.n2139 dvss.t254 28.1205
R6275 dvss.n2103 dvss.t384 28.1205
R6276 dvss.n2067 dvss.t293 28.1205
R6277 dvss.n2031 dvss.t455 28.1205
R6278 dvss.n1998 dvss.t435 28.1205
R6279 dvss.n3367 dvss.t365 28.1205
R6280 dvss.n3270 dvss.t3 28.1205
R6281 dvss.n3155 dvss.t1 28.1205
R6282 dvss.n3041 dvss.t51 28.1205
R6283 dvss.n2922 dvss.t85 28.1205
R6284 dvss.n1427 dvss.t307 28.1205
R6285 dvss.n1330 dvss.t249 28.1205
R6286 dvss.n1053 dvss.t237 28.1205
R6287 dvss.n950 dvss.t194 28.1205
R6288 dvss.n3461 dvss.n3460 27.2737
R6289 dvss.n3312 dvss.n3311 27.2737
R6290 dvss.n3196 dvss.n3195 27.2737
R6291 dvss.n3080 dvss.n3079 27.2737
R6292 dvss.n2964 dvss.n2963 27.2737
R6293 dvss.n1509 dvss.n1470 27.2737
R6294 dvss.n1372 dvss.n1371 27.2737
R6295 dvss.n673 dvss.n672 27.2737
R6296 dvss.n987 dvss.n986 27.2737
R6297 dvss.n2 dvss.t349 24.9236
R6298 dvss.n2 dvss.t500 24.9236
R6299 dvss.n23 dvss.t160 24.9236
R6300 dvss.n23 dvss.t172 24.9236
R6301 dvss.n22 dvss.t152 24.9236
R6302 dvss.n22 dvss.t176 24.9236
R6303 dvss.n30 dvss.t164 24.9236
R6304 dvss.n30 dvss.t166 24.9236
R6305 dvss.n19 dvss.t156 24.9236
R6306 dvss.n19 dvss.t162 24.9236
R6307 dvss.n39 dvss.t148 24.9236
R6308 dvss.n39 dvss.t170 24.9236
R6309 dvss.n16 dvss.t150 24.9236
R6310 dvss.n16 dvss.t174 24.9236
R6311 dvss.n45 dvss.t154 24.9236
R6312 dvss.n45 dvss.t168 24.9236
R6313 dvss.n1980 dvss.n1978 22.5639
R6314 dvss.n3447 dvss.t52 22.5415
R6315 dvss.t26 dvss.n3286 22.5415
R6316 dvss.n3168 dvss.t14 22.5415
R6317 dvss.t4 dvss.n3051 22.5415
R6318 dvss.t278 dvss.n2929 22.5415
R6319 dvss.t372 dvss.n1494 22.5415
R6320 dvss.t469 dvss.n1337 22.5415
R6321 dvss.n1061 dvss.t246 22.5415
R6322 dvss.n857 dvss.t72 22.5415
R6323 dvss.n933 dvss.t256 22.0013
R6324 dvss.n3505 dvss.n3504 21.8222
R6325 dvss.n3331 dvss.n3330 21.8222
R6326 dvss.n3220 dvss.n3219 21.8222
R6327 dvss.n3104 dvss.n3103 21.8222
R6328 dvss.n2983 dvss.n2982 21.8222
R6329 dvss.n1539 dvss.n1538 21.8222
R6330 dvss.n1391 dvss.n1390 21.8222
R6331 dvss.n702 dvss.n701 21.8222
R6332 dvss.n1014 dvss.n1013 21.8222
R6333 dvss.n3618 dvss.n3617 21.8222
R6334 dvss.n2689 dvss.n2688 21.8222
R6335 dvss.n2739 dvss.n2738 21.8222
R6336 dvss.n2789 dvss.n2788 21.8222
R6337 dvss.n2839 dvss.n2838 21.8222
R6338 dvss.n1644 dvss.n1643 21.8222
R6339 dvss.n1249 dvss.n1248 21.8222
R6340 dvss.n1171 dvss.n1170 21.8222
R6341 dvss.n815 dvss.n811 21.8222
R6342 dvss.n93 dvss.t110 21.2805
R6343 dvss.n2293 dvss.t63 21.2805
R6344 dvss.n2207 dvss.t180 21.2805
R6345 dvss.n2175 dvss.t282 21.2805
R6346 dvss.n2139 dvss.t431 21.2805
R6347 dvss.n2103 dvss.t385 21.2805
R6348 dvss.n2067 dvss.t75 21.2805
R6349 dvss.n2031 dvss.t458 21.2805
R6350 dvss.n1998 dvss.t434 21.2805
R6351 dvss.n1979 dvss.t315 21.2805
R6352 dvss.n1979 dvss.t314 21.2805
R6353 dvss.n3367 dvss.t253 21.2805
R6354 dvss.n3270 dvss.t472 21.2805
R6355 dvss.n3155 dvss.t543 21.2805
R6356 dvss.n3041 dvss.t47 21.2805
R6357 dvss.n2922 dvss.t124 21.2805
R6358 dvss.n1427 dvss.t271 21.2805
R6359 dvss.n1330 dvss.t122 21.2805
R6360 dvss.n1053 dvss.t49 21.2805
R6361 dvss.n950 dvss.t460 21.2805
R6362 dvss.n1987 dvss.t309 20.3576
R6363 dvss.n2668 dvss.t495 20.1181
R6364 dvss.n3398 dvss.t104 20.0005
R6365 dvss.n3398 dvss.t108 20.0005
R6366 dvss.n3328 dvss.t490 20.0005
R6367 dvss.n3328 dvss.t452 20.0005
R6368 dvss.n3217 dvss.t140 20.0005
R6369 dvss.n3217 dvss.t454 20.0005
R6370 dvss.n3101 dvss.t537 20.0005
R6371 dvss.n3101 dvss.t413 20.0005
R6372 dvss.n2980 dvss.t209 20.0005
R6373 dvss.n2980 dvss.t514 20.0005
R6374 dvss.n1461 dvss.t264 20.0005
R6375 dvss.n1461 dvss.t319 20.0005
R6376 dvss.n1388 dvss.t518 20.0005
R6377 dvss.n1388 dvss.t439 20.0005
R6378 dvss.n663 dvss.t87 20.0005
R6379 dvss.n663 dvss.t106 20.0005
R6380 dvss.n1011 dvss.t77 20.0005
R6381 dvss.n1011 dvss.t437 20.0005
R6382 dvss.n3612 dvss.t305 20.0005
R6383 dvss.n3612 dvss.t206 20.0005
R6384 dvss.n1773 dvss.t504 20.0005
R6385 dvss.n1773 dvss.t383 20.0005
R6386 dvss.n1742 dvss.t229 20.0005
R6387 dvss.n1742 dvss.t377 20.0005
R6388 dvss.n1711 dvss.t395 20.0005
R6389 dvss.n1711 dvss.t379 20.0005
R6390 dvss.n1680 dvss.t184 20.0005
R6391 dvss.n1680 dvss.t25 20.0005
R6392 dvss.n471 dvss.t333 20.0005
R6393 dvss.n471 dvss.t363 20.0005
R6394 dvss.n1207 dvss.t405 20.0005
R6395 dvss.n1207 dvss.t415 20.0005
R6396 dvss.n581 dvss.t417 20.0005
R6397 dvss.n581 dvss.t251 20.0005
R6398 dvss.n812 dvss.t321 20.0005
R6399 dvss.n812 dvss.t474 20.0005
R6400 dvss.n859 dvss.n856 18.9764
R6401 dvss.n3439 dvss.n3438 18.8324
R6402 dvss.n269 dvss.n259 18.8324
R6403 dvss.n333 dvss.n323 18.8324
R6404 dvss.n3021 dvss.n391 18.8324
R6405 dvss.n2915 dvss.n447 18.8324
R6406 dvss.n1477 dvss.n1476 18.8324
R6407 dvss.n1323 dvss.n556 18.8324
R6408 dvss.n1099 dvss.n626 18.8324
R6409 dvss.n147 dvss.t481 18.3666
R6410 dvss.n1857 dvss.t446 18.3666
R6411 dvss.n2672 dvss.t528 18.3666
R6412 dvss.n1832 dvss.t358 18.3666
R6413 dvss.n1807 dvss.t285 18.3666
R6414 dvss.n1623 dvss.t203 18.3666
R6415 dvss.n1227 dvss.t214 18.3666
R6416 dvss.n1150 dvss.t133 18.3666
R6417 dvss.t44 dvss.n840 18.3666
R6418 dvss.n1048 dvss 18.0711
R6419 dvss dvss.n712 18.0711
R6420 dvss.n1316 dvss 18.0711
R6421 dvss dvss.n554 18.0711
R6422 dvss.n1571 dvss 18.0711
R6423 dvss dvss.n1570 18.0711
R6424 dvss.n2898 dvss 18.0711
R6425 dvss dvss.n445 18.0711
R6426 dvss.n3029 dvss 18.0711
R6427 dvss.n3026 dvss 18.0711
R6428 dvss.n327 dvss 18.0711
R6429 dvss dvss.n321 18.0711
R6430 dvss.n263 dvss 18.0711
R6431 dvss dvss.n257 18.0711
R6432 dvss.n3537 dvss 18.0711
R6433 dvss dvss.n3536 18.0711
R6434 dvss.n3647 dvss 18.0711
R6435 dvss.n2633 dvss 18.0711
R6436 dvss.n2630 dvss 18.0711
R6437 dvss.n2584 dvss 18.0711
R6438 dvss dvss.n2583 18.0711
R6439 dvss.n2537 dvss 18.0711
R6440 dvss dvss.n2536 18.0711
R6441 dvss.n2490 dvss 18.0711
R6442 dvss dvss.n2489 18.0711
R6443 dvss.n2443 dvss 18.0711
R6444 dvss dvss.n2442 18.0711
R6445 dvss.n2396 dvss 18.0711
R6446 dvss dvss.n2395 18.0711
R6447 dvss.n2349 dvss 18.0711
R6448 dvss dvss.n2348 18.0711
R6449 dvss.n2302 dvss 18.0711
R6450 dvss dvss.n2301 18.0711
R6451 dvss.n3700 dvss 18.0711
R6452 dvss dvss.n3699 18.0711
R6453 dvss.n3653 dvss 18.0711
R6454 dvss.n6 dvss.t381 17.4005
R6455 dvss.n6 dvss.t430 17.4005
R6456 dvss.n5 dvss.t345 17.4005
R6457 dvss.n5 dvss.t114 17.4005
R6458 dvss.n1084 dvss.n645 16.2675
R6459 dvss.n3459 dvss.n3423 16.2668
R6460 dvss.n3310 dvss.n238 16.2668
R6461 dvss.n3194 dvss.n3193 16.2668
R6462 dvss.n3078 dvss.n369 16.2668
R6463 dvss.n2962 dvss.n2961 16.2668
R6464 dvss.n1506 dvss.n1505 16.2668
R6465 dvss.n1370 dvss.n1369 16.2668
R6466 dvss.n990 dvss.n748 16.2668
R6467 dvss.n32 dvss.n29 16.132
R6468 dvss.n36 dvss.n20 16.132
R6469 dvss.n41 dvss.n38 16.132
R6470 dvss.n50 dvss.n49 16.132
R6471 dvss.n3750 dvss.n1 16.132
R6472 dvss.n3748 dvss.n3747 16.132
R6473 dvss.n3747 dvss.n3 16.132
R6474 dvss.n27 dvss.n24 15.9567
R6475 dvss.n902 dvss.n901 15.6802
R6476 dvss.n52 dvss.n51 15.606
R6477 dvss.n3743 dvss.n3 15.08
R6478 dvss.n3749 dvss.n3748 14.7293
R6479 dvss.t310 dvss.n902 14.6135
R6480 dvss.n56 dvss.n55 14.5539
R6481 dvss.n52 dvss.n17 13.8526
R6482 dvss.n49 dvss.n46 13.8526
R6483 dvss.n2667 dvss.n2666 13.5291
R6484 dvss.n28 dvss.n27 13.5019
R6485 dvss.n3574 dvss.t485 13.1192
R6486 dvss.t440 dvss.n1851 13.1192
R6487 dvss.t522 dvss.n1881 13.1192
R6488 dvss.t352 dvss.n1826 13.1192
R6489 dvss.n1798 dvss.t289 13.1192
R6490 dvss.t201 dvss.n1606 13.1192
R6491 dvss.n1218 dvss.t220 13.1192
R6492 dvss.t129 dvss.n1133 13.1192
R6493 dvss.n849 dvss.t42 13.1192
R6494 dvss.n3504 dvss.n3397 12.5222
R6495 dvss.n3330 dvss.n3327 12.5222
R6496 dvss.n3219 dvss.n3216 12.5222
R6497 dvss.n3103 dvss.n3100 12.5222
R6498 dvss.n2982 dvss.n2979 12.5222
R6499 dvss.n1538 dvss.n1460 12.5222
R6500 dvss.n1390 dvss.n1387 12.5222
R6501 dvss.n701 dvss.n662 12.5222
R6502 dvss.n1013 dvss.n1010 12.5222
R6503 dvss.n3617 dvss.n3611 12.5222
R6504 dvss.n2688 dvss.n1772 12.5222
R6505 dvss.n2738 dvss.n1741 12.5222
R6506 dvss.n2788 dvss.n1710 12.5222
R6507 dvss.n2838 dvss.n1679 12.5222
R6508 dvss.n1644 dvss.n474 12.5222
R6509 dvss.n1248 dvss.n1206 12.5222
R6510 dvss.n1171 dvss.n584 12.5222
R6511 dvss.n816 dvss.n815 12.5222
R6512 dvss.n2645 dvss.n1980 12.2361
R6513 dvss.n916 dvss.n915 12.1422
R6514 dvss.n3644 dvss.n130 12.0583
R6515 dvss.t240 dvss.n645 11.3665
R6516 dvss.n3459 dvss.t58 11.3663
R6517 dvss.n3310 dvss.t32 11.3663
R6518 dvss.n3194 dvss.t20 11.3663
R6519 dvss.n3078 dvss.t10 11.3663
R6520 dvss.n2962 dvss.t274 11.3663
R6521 dvss.n1505 dvss.t374 11.3663
R6522 dvss.n1370 dvss.t463 11.3663
R6523 dvss.t64 dvss.n748 11.3663
R6524 dvss.n40 dvss.n15 11.0471
R6525 dvss.t74 dvss.t312 10.9522
R6526 dvss.n32 dvss.n31 10.6964
R6527 dvss.n3677 dvss.t96 10.6405
R6528 dvss.n3677 dvss.t100 10.6405
R6529 dvss.n3669 dvss.t94 10.6405
R6530 dvss.n3669 dvss.t102 10.6405
R6531 dvss.n3724 dvss.t492 10.6405
R6532 dvss.n3724 dvss.t488 10.6405
R6533 dvss.n3716 dvss.t496 10.6405
R6534 dvss.n3716 dvss.t498 10.6405
R6535 dvss.n2326 dvss.t142 10.6405
R6536 dvss.n2326 dvss.t136 10.6405
R6537 dvss.n2318 dvss.t144 10.6405
R6538 dvss.n2318 dvss.t138 10.6405
R6539 dvss.n2373 dvss.t532 10.6405
R6540 dvss.n2373 dvss.t533 10.6405
R6541 dvss.n2365 dvss.t539 10.6405
R6542 dvss.n2365 dvss.t535 10.6405
R6543 dvss.n2420 dvss.t213 10.6405
R6544 dvss.n2420 dvss.t212 10.6405
R6545 dvss.n2412 dvss.t211 10.6405
R6546 dvss.n2412 dvss.t210 10.6405
R6547 dvss.n2467 dvss.t269 10.6405
R6548 dvss.n2467 dvss.t265 10.6405
R6549 dvss.n2459 dvss.t268 10.6405
R6550 dvss.n2459 dvss.t267 10.6405
R6551 dvss.n2514 dvss.t521 10.6405
R6552 dvss.n2514 dvss.t520 10.6405
R6553 dvss.n2506 dvss.t519 10.6405
R6554 dvss.n2506 dvss.t515 10.6405
R6555 dvss.n2561 dvss.t92 10.6405
R6556 dvss.n2561 dvss.t91 10.6405
R6557 dvss.n2553 dvss.t90 10.6405
R6558 dvss.n2553 dvss.t89 10.6405
R6559 dvss.n2608 dvss.t83 10.6405
R6560 dvss.n2608 dvss.t82 10.6405
R6561 dvss.n2600 dvss.t81 10.6405
R6562 dvss.n2600 dvss.t80 10.6405
R6563 dvss.n3379 dvss.t57 10.6405
R6564 dvss.n3379 dvss.t59 10.6405
R6565 dvss.n3377 dvss.t53 10.6405
R6566 dvss.n3377 dvss.t55 10.6405
R6567 dvss.n3297 dvss.t31 10.6405
R6568 dvss.n3297 dvss.t33 10.6405
R6569 dvss.n3277 dvss.t27 10.6405
R6570 dvss.n3277 dvss.t29 10.6405
R6571 dvss.n3182 dvss.t19 10.6405
R6572 dvss.n3182 dvss.t21 10.6405
R6573 dvss.n3159 dvss.t15 10.6405
R6574 dvss.n3159 dvss.t17 10.6405
R6575 dvss.n3063 dvss.t9 10.6405
R6576 dvss.n3063 dvss.t11 10.6405
R6577 dvss.n376 dvss.t5 10.6405
R6578 dvss.n376 dvss.t7 10.6405
R6579 dvss.n2949 dvss.t277 10.6405
R6580 dvss.n2949 dvss.t275 10.6405
R6581 dvss.n2935 dvss.t279 10.6405
R6582 dvss.n2935 dvss.t281 10.6405
R6583 dvss.n1439 dvss.t369 10.6405
R6584 dvss.n1439 dvss.t375 10.6405
R6585 dvss.n1437 dvss.t373 10.6405
R6586 dvss.n1437 dvss.t371 10.6405
R6587 dvss.n1357 dvss.t466 10.6405
R6588 dvss.n1357 dvss.t464 10.6405
R6589 dvss.n1343 dvss.t470 10.6405
R6590 dvss.n1343 dvss.t468 10.6405
R6591 dvss.n1073 dvss.t245 10.6405
R6592 dvss.n1073 dvss.t241 10.6405
R6593 dvss.n710 dvss.t247 10.6405
R6594 dvss.n710 dvss.t243 10.6405
R6595 dvss.n743 dvss.t71 10.6405
R6596 dvss.n743 dvss.t65 10.6405
R6597 dvss.n756 dvss.t73 10.6405
R6598 dvss.n756 dvss.t67 10.6405
R6599 dvss.n3402 dvss.t297 10.6405
R6600 dvss.n3402 dvss.t301 10.6405
R6601 dvss.n3498 dvss.t295 10.6405
R6602 dvss.n3498 dvss.t303 10.6405
R6603 dvss.n215 dvss.t506 10.6405
R6604 dvss.n215 dvss.t502 10.6405
R6605 dvss.n218 dvss.t510 10.6405
R6606 dvss.n218 dvss.t512 10.6405
R6607 dvss.n278 dvss.t231 10.6405
R6608 dvss.n278 dvss.t225 10.6405
R6609 dvss.n281 dvss.t233 10.6405
R6610 dvss.n281 dvss.t227 10.6405
R6611 dvss.n342 dvss.t389 10.6405
R6612 dvss.n342 dvss.t391 10.6405
R6613 dvss.n345 dvss.t397 10.6405
R6614 dvss.n345 dvss.t393 10.6405
R6615 dvss.n405 dvss.t192 10.6405
R6616 dvss.n405 dvss.t190 10.6405
R6617 dvss.n408 dvss.t188 10.6405
R6618 dvss.n408 dvss.t186 10.6405
R6619 dvss.n1455 dvss.t343 10.6405
R6620 dvss.n1455 dvss.t335 10.6405
R6621 dvss.n1532 dvss.t341 10.6405
R6622 dvss.n1532 dvss.t339 10.6405
R6623 dvss.n514 dvss.t411 10.6405
R6624 dvss.n514 dvss.t409 10.6405
R6625 dvss.n517 dvss.t407 10.6405
R6626 dvss.n517 dvss.t401 10.6405
R6627 dvss.n657 dvss.t427 10.6405
R6628 dvss.n657 dvss.t425 10.6405
R6629 dvss.n695 dvss.t423 10.6405
R6630 dvss.n695 dvss.t421 10.6405
R6631 dvss.n720 dvss.t331 10.6405
R6632 dvss.n720 dvss.t329 10.6405
R6633 dvss.n723 dvss.t327 10.6405
R6634 dvss.n723 dvss.t325 10.6405
R6635 dvss.n152 dvss.t480 10.6405
R6636 dvss.n152 dvss.t482 10.6405
R6637 dvss.n158 dvss.t486 10.6405
R6638 dvss.n158 dvss.t478 10.6405
R6639 dvss.n1763 dvss.t527 10.6405
R6640 dvss.n1763 dvss.t529 10.6405
R6641 dvss.n1757 dvss.t523 10.6405
R6642 dvss.n1757 dvss.t525 10.6405
R6643 dvss.n1732 dvss.t445 10.6405
R6644 dvss.n1732 dvss.t447 10.6405
R6645 dvss.n1726 dvss.t441 10.6405
R6646 dvss.n1726 dvss.t443 10.6405
R6647 dvss.n1701 dvss.t357 10.6405
R6648 dvss.n1701 dvss.t359 10.6405
R6649 dvss.n1695 dvss.t353 10.6405
R6650 dvss.n1695 dvss.t355 10.6405
R6651 dvss.n1670 dvss.t288 10.6405
R6652 dvss.n1670 dvss.t286 10.6405
R6653 dvss.n1663 dvss.t290 10.6405
R6654 dvss.n1663 dvss.t292 10.6405
R6655 dvss.n481 dvss.t198 10.6405
R6656 dvss.n481 dvss.t204 10.6405
R6657 dvss.n490 dvss.t202 10.6405
R6658 dvss.n490 dvss.t200 10.6405
R6659 dvss.n1197 dvss.t217 10.6405
R6660 dvss.n1197 dvss.t215 10.6405
R6661 dvss.n1190 dvss.t221 10.6405
R6662 dvss.n1190 dvss.t219 10.6405
R6663 dvss.n591 dvss.t128 10.6405
R6664 dvss.n591 dvss.t134 10.6405
R6665 dvss.n600 dvss.t130 10.6405
R6666 dvss.n600 dvss.t126 10.6405
R6667 dvss.n794 dvss.t41 10.6405
R6668 dvss.n794 dvss.t45 10.6405
R6669 dvss.n784 dvss.t43 10.6405
R6670 dvss.n784 dvss.t37 10.6405
R6671 dvss.n3378 dvss.n3376 10.64
R6672 dvss.n3282 dvss.n3281 10.64
R6673 dvss.n3164 dvss.n3163 10.64
R6674 dvss.n385 dvss.n377 10.64
R6675 dvss.n2936 dvss.n2934 10.64
R6676 dvss.n1438 dvss.n1436 10.64
R6677 dvss.n1344 dvss.n1342 10.64
R6678 dvss.n711 dvss.n709 10.64
R6679 dvss.n964 dvss.n757 10.64
R6680 dvss.n3578 dvss.n159 10.64
R6681 dvss.n2715 dvss.n2714 10.64
R6682 dvss.n2765 dvss.n2764 10.64
R6683 dvss.n2815 dvss.n2814 10.64
R6684 dvss.n2865 dvss.n2864 10.64
R6685 dvss.n1600 dvss.n491 10.64
R6686 dvss.n1275 dvss.n1274 10.64
R6687 dvss.n1127 dvss.n601 10.64
R6688 dvss.n787 dvss.n785 10.64
R6689 dvss.t312 dvss.t308 10.6301
R6690 dvss.n3744 dvss.n3743 10.3526
R6691 dvss.n898 dvss 9.3467
R6692 dvss.n2664 dvss 9.3467
R6693 dvss.n814 dvss.n813 9.3005
R6694 dvss.n817 dvss.n816 9.3005
R6695 dvss.n801 dvss.n800 9.3005
R6696 dvss.n790 dvss.n789 9.3005
R6697 dvss.n793 dvss.n792 9.3005
R6698 dvss.n798 dvss.n797 9.3005
R6699 dvss.n802 dvss.n801 9.3005
R6700 dvss.n1173 dvss.n1172 9.3005
R6701 dvss.n584 dvss.n583 9.3005
R6702 dvss.n1157 dvss.n589 9.3005
R6703 dvss.n1140 dvss.n1139 9.3005
R6704 dvss.n1143 dvss.n1142 9.3005
R6705 dvss.n1155 dvss.n1154 9.3005
R6706 dvss.n1158 dvss.n1157 9.3005
R6707 dvss.n1247 dvss.n1246 9.3005
R6708 dvss.n1245 dvss.n1206 9.3005
R6709 dvss.n1258 dvss.n1257 9.3005
R6710 dvss.n1273 dvss.n1272 9.3005
R6711 dvss.n1267 dvss.n1266 9.3005
R6712 dvss.n1264 dvss.n1263 9.3005
R6713 dvss.n1257 dvss.n1255 9.3005
R6714 dvss.n1646 dvss.n1645 9.3005
R6715 dvss.n474 dvss.n473 9.3005
R6716 dvss.n1630 dvss.n479 9.3005
R6717 dvss.n1613 dvss.n1612 9.3005
R6718 dvss.n1616 dvss.n1615 9.3005
R6719 dvss.n1628 dvss.n1627 9.3005
R6720 dvss.n1631 dvss.n1630 9.3005
R6721 dvss.n2837 dvss.n2836 9.3005
R6722 dvss.n2835 dvss.n1679 9.3005
R6723 dvss.n2848 dvss.n2847 9.3005
R6724 dvss.n2863 dvss.n2862 9.3005
R6725 dvss.n2857 dvss.n2856 9.3005
R6726 dvss.n2854 dvss.n2853 9.3005
R6727 dvss.n2847 dvss.n2845 9.3005
R6728 dvss.n2787 dvss.n2786 9.3005
R6729 dvss.n2785 dvss.n1710 9.3005
R6730 dvss.n2798 dvss.n2797 9.3005
R6731 dvss.n2813 dvss.n2812 9.3005
R6732 dvss.n2807 dvss.n2806 9.3005
R6733 dvss.n2804 dvss.n2803 9.3005
R6734 dvss.n2797 dvss.n2795 9.3005
R6735 dvss.n2737 dvss.n2736 9.3005
R6736 dvss.n2735 dvss.n1741 9.3005
R6737 dvss.n2748 dvss.n2747 9.3005
R6738 dvss.n2763 dvss.n2762 9.3005
R6739 dvss.n2757 dvss.n2756 9.3005
R6740 dvss.n2754 dvss.n2753 9.3005
R6741 dvss.n2747 dvss.n2745 9.3005
R6742 dvss.n2687 dvss.n2686 9.3005
R6743 dvss.n2685 dvss.n1772 9.3005
R6744 dvss.n2698 dvss.n2697 9.3005
R6745 dvss.n2713 dvss.n2712 9.3005
R6746 dvss.n2707 dvss.n2706 9.3005
R6747 dvss.n2704 dvss.n2703 9.3005
R6748 dvss.n2697 dvss.n2695 9.3005
R6749 dvss.n3616 dvss.n3615 9.3005
R6750 dvss.n3614 dvss.n3611 9.3005
R6751 dvss.n3600 dvss.n3599 9.3005
R6752 dvss.n3581 dvss.n3580 9.3005
R6753 dvss.n3584 dvss.n3583 9.3005
R6754 dvss.n3597 dvss.n3596 9.3005
R6755 dvss.n3599 dvss.n151 9.3005
R6756 dvss.n953 dvss.n952 9.3005
R6757 dvss.n954 dvss.n953 9.3005
R6758 dvss.n1038 dvss.n1037 9.3005
R6759 dvss.n1039 dvss.n1038 9.3005
R6760 dvss.n1035 dvss.n722 9.3005
R6761 dvss.n1035 dvss.n1034 9.3005
R6762 dvss.n737 dvss.n721 9.3005
R6763 dvss.n999 dvss.n721 9.3005
R6764 dvss.n1056 dvss.n1055 9.3005
R6765 dvss.n1057 dvss.n1056 9.3005
R6766 dvss.n1299 dvss.n1298 9.3005
R6767 dvss.n1298 dvss.n1297 9.3005
R6768 dvss.n698 dvss.n697 9.3005
R6769 dvss.n697 dvss.n696 9.3005
R6770 dvss.n659 dvss.n658 9.3005
R6771 dvss.n658 dvss.n652 9.3005
R6772 dvss.n1333 dvss.n1332 9.3005
R6773 dvss.n1332 dvss.n1329 9.3005
R6774 dvss.n1414 dvss.n511 9.3005
R6775 dvss.n1415 dvss.n1414 9.3005
R6776 dvss.n1412 dvss.n516 9.3005
R6777 dvss.n1412 dvss.n1411 9.3005
R6778 dvss.n1382 dvss.n515 9.3005
R6779 dvss.n532 dvss.n515 9.3005
R6780 dvss.n1566 dvss.n1565 9.3005
R6781 dvss.n1567 dvss.n1566 9.3005
R6782 dvss.n2889 dvss.n2888 9.3005
R6783 dvss.n2888 dvss.n2887 9.3005
R6784 dvss.n1535 dvss.n1534 9.3005
R6785 dvss.n1534 dvss.n1533 9.3005
R6786 dvss.n1457 dvss.n1456 9.3005
R6787 dvss.n1456 dvss.n1449 9.3005
R6788 dvss.n2925 dvss.n2924 9.3005
R6789 dvss.n2924 dvss.n2921 9.3005
R6790 dvss.n3007 dvss.n401 9.3005
R6791 dvss.n3008 dvss.n3007 9.3005
R6792 dvss.n3005 dvss.n407 9.3005
R6793 dvss.n3005 dvss.n3004 9.3005
R6794 dvss.n2974 dvss.n406 9.3005
R6795 dvss.n423 dvss.n406 9.3005
R6796 dvss.n3044 dvss.n3043 9.3005
R6797 dvss.n3043 dvss.n3040 9.3005
R6798 dvss.n3124 dvss.n339 9.3005
R6799 dvss.n3125 dvss.n3124 9.3005
R6800 dvss.n3122 dvss.n344 9.3005
R6801 dvss.n3122 dvss.n3121 9.3005
R6802 dvss.n3090 dvss.n343 9.3005
R6803 dvss.n363 dvss.n343 9.3005
R6804 dvss.n3158 dvss.n3157 9.3005
R6805 dvss.n3157 dvss.n3154 9.3005
R6806 dvss.n3240 dvss.n275 9.3005
R6807 dvss.n3241 dvss.n3240 9.3005
R6808 dvss.n3238 dvss.n280 9.3005
R6809 dvss.n3238 dvss.n3237 9.3005
R6810 dvss.n3206 dvss.n279 9.3005
R6811 dvss.n299 dvss.n279 9.3005
R6812 dvss.n3273 dvss.n3272 9.3005
R6813 dvss.n3272 dvss.n3269 9.3005
R6814 dvss.n3354 dvss.n212 9.3005
R6815 dvss.n3355 dvss.n3354 9.3005
R6816 dvss.n3352 dvss.n217 9.3005
R6817 dvss.n3352 dvss.n3351 9.3005
R6818 dvss.n3322 dvss.n216 9.3005
R6819 dvss.n233 dvss.n216 9.3005
R6820 dvss.n3532 dvss.n3531 9.3005
R6821 dvss.n3533 dvss.n3532 9.3005
R6822 dvss.n3496 dvss.n3495 9.3005
R6823 dvss.n3496 dvss.n3404 9.3005
R6824 dvss.n3501 dvss.n3500 9.3005
R6825 dvss.n3500 dvss.n3499 9.3005
R6826 dvss.n3403 dvss.n3401 9.3005
R6827 dvss.n3403 dvss.n3389 9.3005
R6828 dvss.n912 dvss.n911 9.3005
R6829 dvss.n911 dvss.n910 9.3005
R6830 dvss.n936 dvss.n935 9.3005
R6831 dvss.n935 dvss.n934 9.3005
R6832 dvss.n1012 dvss.n725 9.3005
R6833 dvss.n1010 dvss.n1009 9.3005
R6834 dvss.n997 dvss.n742 9.3005
R6835 dvss.n974 dvss.n973 9.3005
R6836 dvss.n977 dvss.n976 9.3005
R6837 dvss.n995 dvss.n994 9.3005
R6838 dvss.n998 dvss.n997 9.3005
R6839 dvss.n700 dvss.n699 9.3005
R6840 dvss.n694 dvss.n662 9.3005
R6841 dvss.n1079 dvss.n1078 9.3005
R6842 dvss.n1069 dvss.n1068 9.3005
R6843 dvss.n1072 dvss.n1071 9.3005
R6844 dvss.n1076 dvss.n1075 9.3005
R6845 dvss.n1078 dvss.n708 9.3005
R6846 dvss.n1389 dvss.n519 9.3005
R6847 dvss.n1387 dvss.n1386 9.3005
R6848 dvss.n1380 dvss.n1379 9.3005
R6849 dvss.n1346 dvss.n1345 9.3005
R6850 dvss.n1356 dvss.n1355 9.3005
R6851 dvss.n1361 dvss.n1360 9.3005
R6852 dvss.n1381 dvss.n1380 9.3005
R6853 dvss.n1537 dvss.n1536 9.3005
R6854 dvss.n1531 dvss.n1460 9.3005
R6855 dvss.n1550 dvss.n1549 9.3005
R6856 dvss.n1560 dvss.n1559 9.3005
R6857 dvss.n1557 dvss.n1556 9.3005
R6858 dvss.n1547 dvss.n1546 9.3005
R6859 dvss.n1549 dvss.n1545 9.3005
R6860 dvss.n2981 dvss.n410 9.3005
R6861 dvss.n2979 dvss.n2978 9.3005
R6862 dvss.n2972 dvss.n2971 9.3005
R6863 dvss.n2938 dvss.n2937 9.3005
R6864 dvss.n2948 dvss.n2947 9.3005
R6865 dvss.n2953 dvss.n2952 9.3005
R6866 dvss.n2973 dvss.n2972 9.3005
R6867 dvss.n3102 dvss.n347 9.3005
R6868 dvss.n3100 dvss.n3099 9.3005
R6869 dvss.n3088 dvss.n3087 9.3005
R6870 dvss.n3061 dvss.n3060 9.3005
R6871 dvss.n3070 dvss.n3069 9.3005
R6872 dvss.n3067 dvss.n3066 9.3005
R6873 dvss.n3089 dvss.n3088 9.3005
R6874 dvss.n3218 dvss.n283 9.3005
R6875 dvss.n3216 dvss.n3215 9.3005
R6876 dvss.n3204 dvss.n3203 9.3005
R6877 dvss.n3162 dvss.n3161 9.3005
R6878 dvss.n3181 dvss.n3180 9.3005
R6879 dvss.n3186 dvss.n3185 9.3005
R6880 dvss.n3205 dvss.n3204 9.3005
R6881 dvss.n3329 dvss.n220 9.3005
R6882 dvss.n3327 dvss.n3326 9.3005
R6883 dvss.n3320 dvss.n3319 9.3005
R6884 dvss.n3280 dvss.n3279 9.3005
R6885 dvss.n3296 dvss.n3295 9.3005
R6886 dvss.n3301 dvss.n3300 9.3005
R6887 dvss.n3321 dvss.n3320 9.3005
R6888 dvss.n3503 dvss.n3502 9.3005
R6889 dvss.n3400 dvss.n3397 9.3005
R6890 dvss.n3516 dvss.n3515 9.3005
R6891 dvss.n3526 dvss.n3525 9.3005
R6892 dvss.n3523 dvss.n3522 9.3005
R6893 dvss.n3513 dvss.n3512 9.3005
R6894 dvss.n3515 dvss.n3511 9.3005
R6895 dvss.n916 dvss.n868 9.3005
R6896 dvss.n917 dvss.n916 9.3005
R6897 dvss.n897 dvss.n878 9.3005
R6898 dvss.n896 dvss.n879 9.3005
R6899 dvss.n884 dvss.n880 9.3005
R6900 dvss.n890 dvss.n886 9.3005
R6901 dvss.n889 dvss.n888 9.3005
R6902 dvss.n887 dvss.n873 9.3005
R6903 dvss.n909 dvss.n908 9.3005
R6904 dvss.n913 dvss.n872 9.3005
R6905 dvss.n920 dvss.n919 9.3005
R6906 dvss.n918 dvss.n869 9.3005
R6907 dvss.n928 dvss.n927 9.3005
R6908 dvss.n929 dvss.n867 9.3005
R6909 dvss.n939 dvss.n930 9.3005
R6910 dvss.n938 dvss.n937 9.3005
R6911 dvss.n932 dvss.n865 9.3005
R6912 dvss.n931 dvss.n862 9.3005
R6913 dvss.n949 dvss.n948 9.3005
R6914 dvss.n955 dvss.n762 9.3005
R6915 dvss.n961 dvss.n763 9.3005
R6916 dvss.n963 dvss.n962 9.3005
R6917 dvss.n965 dvss.n758 9.3005
R6918 dvss.n972 dvss.n971 9.3005
R6919 dvss.n978 dvss.n754 9.3005
R6920 dvss.n755 dvss.n750 9.3005
R6921 dvss.n993 dvss.n745 9.3005
R6922 dvss.n985 dvss.n984 9.3005
R6923 dvss.n1000 dvss.n736 9.3005
R6924 dvss.n1007 dvss.n738 9.3005
R6925 dvss.n1016 dvss.n1008 9.3005
R6926 dvss.n1015 dvss.n732 9.3005
R6927 dvss.n1033 dvss.n724 9.3005
R6928 dvss.n1030 dvss.n729 9.3005
R6929 dvss.n1029 dvss.n1028 9.3005
R6930 dvss.n1040 dvss.n619 9.3005
R6931 dvss.n1105 dvss.n620 9.3005
R6932 dvss.n1104 dvss.n621 9.3005
R6933 dvss.n1103 dvss.n622 9.3005
R6934 dvss.n1049 dvss.n623 9.3005
R6935 dvss.n1052 dvss.n1051 9.3005
R6936 dvss.n1058 dvss.n630 9.3005
R6937 dvss.n1096 dvss.n631 9.3005
R6938 dvss.n1095 dvss.n632 9.3005
R6939 dvss.n1094 dvss.n633 9.3005
R6940 dvss.n1067 dvss.n634 9.3005
R6941 dvss.n1088 dvss.n640 9.3005
R6942 dvss.n1087 dvss.n641 9.3005
R6943 dvss.n1086 dvss.n642 9.3005
R6944 dvss.n1080 dvss.n643 9.3005
R6945 dvss.n670 dvss.n651 9.3005
R6946 dvss.n707 dvss.n653 9.3005
R6947 dvss.n704 dvss.n660 9.3005
R6948 dvss.n703 dvss.n661 9.3005
R6949 dvss.n669 dvss.n664 9.3005
R6950 dvss.n693 dvss.n665 9.3005
R6951 dvss.n690 dvss.n568 9.3005
R6952 dvss.n1296 dvss.n1295 9.3005
R6953 dvss.n1300 dvss.n562 9.3005
R6954 dvss.n1320 dvss.n563 9.3005
R6955 dvss.n1319 dvss.n1318 9.3005
R6956 dvss.n1315 dvss.n564 9.3005
R6957 dvss.n1314 dvss.n1313 9.3005
R6958 dvss.n1328 dvss.n553 9.3005
R6959 dvss.n552 dvss.n551 9.3005
R6960 dvss.n1335 dvss.n1334 9.3005
R6961 dvss.n1341 dvss.n547 9.3005
R6962 dvss.n1348 dvss.n1347 9.3005
R6963 dvss.n1354 dvss.n539 9.3005
R6964 dvss.n1363 dvss.n1362 9.3005
R6965 dvss.n1366 dvss.n1364 9.3005
R6966 dvss.n1365 dvss.n536 9.3005
R6967 dvss.n1378 dvss.n530 9.3005
R6968 dvss.n1384 dvss.n1383 9.3005
R6969 dvss.n1393 dvss.n1385 9.3005
R6970 dvss.n1392 dvss.n526 9.3005
R6971 dvss.n1410 dvss.n518 9.3005
R6972 dvss.n1407 dvss.n523 9.3005
R6973 dvss.n1406 dvss.n1405 9.3005
R6974 dvss.n1416 dvss.n509 9.3005
R6975 dvss.n1578 dvss.n1577 9.3005
R6976 dvss.n1574 dvss.n510 9.3005
R6977 dvss.n1573 dvss.n1420 9.3005
R6978 dvss.n1572 dvss.n1421 9.3005
R6979 dvss.n1569 dvss.n1425 9.3005
R6980 dvss.n1568 dvss.n1426 9.3005
R6981 dvss.n1491 dvss.n1429 9.3005
R6982 dvss.n1564 dvss.n1430 9.3005
R6983 dvss.n1561 dvss.n1435 9.3005
R6984 dvss.n1499 dvss.n1498 9.3005
R6985 dvss.n1501 dvss.n1500 9.3005
R6986 dvss.n1555 dvss.n1441 9.3005
R6987 dvss.n1552 dvss.n1446 9.3005
R6988 dvss.n1551 dvss.n1447 9.3005
R6989 dvss.n1468 dvss.n1448 9.3005
R6990 dvss.n1544 dvss.n1450 9.3005
R6991 dvss.n1541 dvss.n1458 9.3005
R6992 dvss.n1540 dvss.n1459 9.3005
R6993 dvss.n1467 dvss.n1462 9.3005
R6994 dvss.n1530 dvss.n1463 9.3005
R6995 dvss.n1527 dvss.n458 9.3005
R6996 dvss.n2886 dvss.n2885 9.3005
R6997 dvss.n2890 dvss.n453 9.3005
R6998 dvss.n2912 dvss.n2911 9.3005
R6999 dvss.n2908 dvss.n454 9.3005
R7000 dvss.n2907 dvss.n2899 9.3005
R7001 dvss.n2906 dvss.n2905 9.3005
R7002 dvss.n2920 dvss.n444 9.3005
R7003 dvss.n443 dvss.n442 9.3005
R7004 dvss.n2927 dvss.n2926 9.3005
R7005 dvss.n2933 dvss.n438 9.3005
R7006 dvss.n2940 dvss.n2939 9.3005
R7007 dvss.n2946 dvss.n430 9.3005
R7008 dvss.n2955 dvss.n2954 9.3005
R7009 dvss.n2958 dvss.n2956 9.3005
R7010 dvss.n2957 dvss.n427 9.3005
R7011 dvss.n2970 dvss.n421 9.3005
R7012 dvss.n2976 dvss.n2975 9.3005
R7013 dvss.n2985 dvss.n2977 9.3005
R7014 dvss.n2984 dvss.n417 9.3005
R7015 dvss.n3003 dvss.n409 9.3005
R7016 dvss.n3000 dvss.n414 9.3005
R7017 dvss.n2999 dvss.n2998 9.3005
R7018 dvss.n3009 dvss.n400 9.3005
R7019 dvss.n3013 dvss.n3012 9.3005
R7020 dvss.n402 dvss.n394 9.3005
R7021 dvss.n3032 dvss.n3031 9.3005
R7022 dvss.n3028 dvss.n395 9.3005
R7023 dvss.n3027 dvss.n388 9.3005
R7024 dvss.n3039 dvss.n3038 9.3005
R7025 dvss.n3045 dvss.n383 9.3005
R7026 dvss.n3049 dvss.n3048 9.3005
R7027 dvss.n384 dvss.n378 9.3005
R7028 dvss.n3059 dvss.n3058 9.3005
R7029 dvss.n3071 dvss.n373 9.3005
R7030 dvss.n3075 dvss.n3074 9.3005
R7031 dvss.n3065 dvss.n366 9.3005
R7032 dvss.n3083 dvss.n3082 9.3005
R7033 dvss.n3086 dvss.n362 9.3005
R7034 dvss.n3092 dvss.n3091 9.3005
R7035 dvss.n3098 dvss.n357 9.3005
R7036 dvss.n3106 dvss.n3105 9.3005
R7037 dvss.n3120 dvss.n346 9.3005
R7038 dvss.n3117 dvss.n3115 9.3005
R7039 dvss.n3116 dvss.n340 9.3005
R7040 dvss.n3127 dvss.n3126 9.3005
R7041 dvss.n3130 dvss.n3128 9.3005
R7042 dvss.n3129 dvss.n335 9.3005
R7043 dvss.n3144 dvss.n328 9.3005
R7044 dvss.n3143 dvss.n329 9.3005
R7045 dvss.n3142 dvss.n3141 9.3005
R7046 dvss.n3153 dvss.n320 9.3005
R7047 dvss.n319 dvss.n318 9.3005
R7048 dvss.n3166 dvss.n3165 9.3005
R7049 dvss.n3160 dvss.n313 9.3005
R7050 dvss.n3176 dvss.n3175 9.3005
R7051 dvss.n3179 dvss.n308 9.3005
R7052 dvss.n3188 dvss.n3187 9.3005
R7053 dvss.n309 dvss.n302 9.3005
R7054 dvss.n3199 dvss.n3198 9.3005
R7055 dvss.n3202 dvss.n298 9.3005
R7056 dvss.n3208 dvss.n3207 9.3005
R7057 dvss.n3214 dvss.n293 9.3005
R7058 dvss.n3222 dvss.n3221 9.3005
R7059 dvss.n3236 dvss.n282 9.3005
R7060 dvss.n3233 dvss.n3231 9.3005
R7061 dvss.n3232 dvss.n276 9.3005
R7062 dvss.n3243 dvss.n3242 9.3005
R7063 dvss.n3246 dvss.n3244 9.3005
R7064 dvss.n3245 dvss.n271 9.3005
R7065 dvss.n3260 dvss.n264 9.3005
R7066 dvss.n3259 dvss.n265 9.3005
R7067 dvss.n3258 dvss.n3257 9.3005
R7068 dvss.n3268 dvss.n255 9.3005
R7069 dvss.n3275 dvss.n3274 9.3005
R7070 dvss.n3283 dvss.n3276 9.3005
R7071 dvss.n3278 dvss.n252 9.3005
R7072 dvss.n3293 dvss.n246 9.3005
R7073 dvss.n3294 dvss.n241 9.3005
R7074 dvss.n3307 dvss.n3306 9.3005
R7075 dvss.n3303 dvss.n242 9.3005
R7076 dvss.n3302 dvss.n237 9.3005
R7077 dvss.n3318 dvss.n231 9.3005
R7078 dvss.n3324 dvss.n3323 9.3005
R7079 dvss.n3333 dvss.n3325 9.3005
R7080 dvss.n3332 dvss.n227 9.3005
R7081 dvss.n3350 dvss.n219 9.3005
R7082 dvss.n3347 dvss.n224 9.3005
R7083 dvss.n3346 dvss.n3345 9.3005
R7084 dvss.n3356 dvss.n210 9.3005
R7085 dvss.n3544 dvss.n3543 9.3005
R7086 dvss.n3540 dvss.n211 9.3005
R7087 dvss.n3539 dvss.n3360 9.3005
R7088 dvss.n3538 dvss.n3361 9.3005
R7089 dvss.n3535 dvss.n3365 9.3005
R7090 dvss.n3534 dvss.n3366 9.3005
R7091 dvss.n3429 dvss.n3369 9.3005
R7092 dvss.n3530 dvss.n3370 9.3005
R7093 dvss.n3527 dvss.n3375 9.3005
R7094 dvss.n3426 dvss.n3425 9.3005
R7095 dvss.n3428 dvss.n3427 9.3005
R7096 dvss.n3521 dvss.n3381 9.3005
R7097 dvss.n3518 dvss.n3386 9.3005
R7098 dvss.n3517 dvss.n3387 9.3005
R7099 dvss.n3422 dvss.n3388 9.3005
R7100 dvss.n3510 dvss.n3390 9.3005
R7101 dvss.n3507 dvss.n3395 9.3005
R7102 dvss.n3506 dvss.n3396 9.3005
R7103 dvss.n3415 dvss.n3399 9.3005
R7104 dvss.n3476 dvss.n3475 9.3005
R7105 dvss.n3418 dvss.n3416 9.3005
R7106 dvss.n3417 dvss.n3411 9.3005
R7107 dvss.n3494 dvss.n3405 9.3005
R7108 dvss.n3491 dvss.n3409 9.3005
R7109 dvss.n3490 dvss.n3489 9.3005
R7110 dvss.n3646 dvss.n125 9.3005
R7111 dvss.n854 dvss.n768 9.3005
R7112 dvss.n853 dvss.n769 9.3005
R7113 dvss.n852 dvss.n770 9.3005
R7114 dvss.n786 dvss.n771 9.3005
R7115 dvss.n788 dvss.n775 9.3005
R7116 dvss.n845 dvss.n776 9.3005
R7117 dvss.n844 dvss.n777 9.3005
R7118 dvss.n843 dvss.n778 9.3005
R7119 dvss.n796 dvss.n779 9.3005
R7120 dvss.n837 dvss.n782 9.3005
R7121 dvss.n836 dvss.n783 9.3005
R7122 dvss.n835 dvss.n803 9.3005
R7123 dvss.n808 dvss.n804 9.3005
R7124 dvss.n829 dvss.n809 9.3005
R7125 dvss.n828 dvss.n810 9.3005
R7126 dvss.n827 dvss.n818 9.3005
R7127 dvss.n821 dvss.n820 9.3005
R7128 dvss.n819 dvss.n611 9.3005
R7129 dvss.n1114 dvss.n1113 9.3005
R7130 dvss.n1115 dvss.n610 9.3005
R7131 dvss.n1118 dvss.n1117 9.3005
R7132 dvss.n1116 dvss.n607 9.3005
R7133 dvss.n1125 dvss.n1124 9.3005
R7134 dvss.n1126 dvss.n606 9.3005
R7135 dvss.n1130 dvss.n1129 9.3005
R7136 dvss.n1128 dvss.n602 9.3005
R7137 dvss.n1137 dvss.n1136 9.3005
R7138 dvss.n1138 dvss.n598 9.3005
R7139 dvss.n1145 dvss.n1144 9.3005
R7140 dvss.n599 dvss.n594 9.3005
R7141 dvss.n1153 dvss.n1152 9.3005
R7142 dvss.n593 dvss.n588 9.3005
R7143 dvss.n1160 dvss.n1159 9.3005
R7144 dvss.n590 dvss.n585 9.3005
R7145 dvss.n1168 dvss.n1167 9.3005
R7146 dvss.n1169 dvss.n580 9.3005
R7147 dvss.n1175 dvss.n1174 9.3005
R7148 dvss.n582 dvss.n577 9.3005
R7149 dvss.n1182 dvss.n1181 9.3005
R7150 dvss.n1183 dvss.n575 9.3005
R7151 dvss.n1288 dvss.n1287 9.3005
R7152 dvss.n1286 dvss.n576 9.3005
R7153 dvss.n1285 dvss.n1284 9.3005
R7154 dvss.n1283 dvss.n1282 9.3005
R7155 dvss.n1281 dvss.n1186 9.3005
R7156 dvss.n1280 dvss.n1279 9.3005
R7157 dvss.n1278 dvss.n1277 9.3005
R7158 dvss.n1276 dvss.n1189 9.3005
R7159 dvss.n1192 dvss.n1191 9.3005
R7160 dvss.n1271 dvss.n1270 9.3005
R7161 dvss.n1269 dvss.n1268 9.3005
R7162 dvss.n1198 dvss.n1195 9.3005
R7163 dvss.n1262 dvss.n1261 9.3005
R7164 dvss.n1260 dvss.n1259 9.3005
R7165 dvss.n1202 dvss.n1201 9.3005
R7166 dvss.n1254 dvss.n1253 9.3005
R7167 dvss.n1252 dvss.n1251 9.3005
R7168 dvss.n1250 dvss.n1205 9.3005
R7169 dvss.n1209 dvss.n1208 9.3005
R7170 dvss.n1244 dvss.n1243 9.3005
R7171 dvss.n1242 dvss.n1241 9.3005
R7172 dvss.n1240 dvss.n501 9.3005
R7173 dvss.n1587 dvss.n1586 9.3005
R7174 dvss.n1588 dvss.n500 9.3005
R7175 dvss.n1591 dvss.n1590 9.3005
R7176 dvss.n1589 dvss.n497 9.3005
R7177 dvss.n1598 dvss.n1597 9.3005
R7178 dvss.n1599 dvss.n496 9.3005
R7179 dvss.n1603 dvss.n1602 9.3005
R7180 dvss.n1601 dvss.n492 9.3005
R7181 dvss.n1610 dvss.n1609 9.3005
R7182 dvss.n1611 dvss.n488 9.3005
R7183 dvss.n1618 dvss.n1617 9.3005
R7184 dvss.n489 dvss.n484 9.3005
R7185 dvss.n1626 dvss.n1625 9.3005
R7186 dvss.n483 dvss.n478 9.3005
R7187 dvss.n1633 dvss.n1632 9.3005
R7188 dvss.n480 dvss.n475 9.3005
R7189 dvss.n1641 dvss.n1640 9.3005
R7190 dvss.n1642 dvss.n470 9.3005
R7191 dvss.n1648 dvss.n1647 9.3005
R7192 dvss.n472 dvss.n467 9.3005
R7193 dvss.n1655 dvss.n1654 9.3005
R7194 dvss.n1656 dvss.n465 9.3005
R7195 dvss.n2878 dvss.n2877 9.3005
R7196 dvss.n2876 dvss.n466 9.3005
R7197 dvss.n2875 dvss.n2874 9.3005
R7198 dvss.n2873 dvss.n2872 9.3005
R7199 dvss.n2871 dvss.n1659 9.3005
R7200 dvss.n2870 dvss.n2869 9.3005
R7201 dvss.n2868 dvss.n2867 9.3005
R7202 dvss.n2866 dvss.n1662 9.3005
R7203 dvss.n1665 dvss.n1664 9.3005
R7204 dvss.n2861 dvss.n2860 9.3005
R7205 dvss.n2859 dvss.n2858 9.3005
R7206 dvss.n1671 dvss.n1668 9.3005
R7207 dvss.n2852 dvss.n2851 9.3005
R7208 dvss.n2850 dvss.n2849 9.3005
R7209 dvss.n1675 dvss.n1674 9.3005
R7210 dvss.n2844 dvss.n2843 9.3005
R7211 dvss.n2842 dvss.n2841 9.3005
R7212 dvss.n2840 dvss.n1678 9.3005
R7213 dvss.n1682 dvss.n1681 9.3005
R7214 dvss.n2834 dvss.n2833 9.3005
R7215 dvss.n2832 dvss.n2831 9.3005
R7216 dvss.n2830 dvss.n1685 9.3005
R7217 dvss.n2829 dvss.n2828 9.3005
R7218 dvss.n2827 dvss.n2826 9.3005
R7219 dvss.n2825 dvss.n1688 9.3005
R7220 dvss.n2824 dvss.n2823 9.3005
R7221 dvss.n2822 dvss.n2821 9.3005
R7222 dvss.n2820 dvss.n1691 9.3005
R7223 dvss.n2819 dvss.n2818 9.3005
R7224 dvss.n2817 dvss.n2816 9.3005
R7225 dvss.n1696 dvss.n1694 9.3005
R7226 dvss.n2811 dvss.n2810 9.3005
R7227 dvss.n2809 dvss.n2808 9.3005
R7228 dvss.n1702 dvss.n1699 9.3005
R7229 dvss.n2802 dvss.n2801 9.3005
R7230 dvss.n2800 dvss.n2799 9.3005
R7231 dvss.n1706 dvss.n1705 9.3005
R7232 dvss.n2794 dvss.n2793 9.3005
R7233 dvss.n2792 dvss.n2791 9.3005
R7234 dvss.n2790 dvss.n1709 9.3005
R7235 dvss.n1713 dvss.n1712 9.3005
R7236 dvss.n2784 dvss.n2783 9.3005
R7237 dvss.n2782 dvss.n2781 9.3005
R7238 dvss.n2780 dvss.n1716 9.3005
R7239 dvss.n2779 dvss.n2778 9.3005
R7240 dvss.n2777 dvss.n2776 9.3005
R7241 dvss.n2775 dvss.n1719 9.3005
R7242 dvss.n2774 dvss.n2773 9.3005
R7243 dvss.n2772 dvss.n2771 9.3005
R7244 dvss.n2770 dvss.n1722 9.3005
R7245 dvss.n2769 dvss.n2768 9.3005
R7246 dvss.n2767 dvss.n2766 9.3005
R7247 dvss.n1727 dvss.n1725 9.3005
R7248 dvss.n2761 dvss.n2760 9.3005
R7249 dvss.n2759 dvss.n2758 9.3005
R7250 dvss.n1733 dvss.n1730 9.3005
R7251 dvss.n2752 dvss.n2751 9.3005
R7252 dvss.n2750 dvss.n2749 9.3005
R7253 dvss.n1737 dvss.n1736 9.3005
R7254 dvss.n2744 dvss.n2743 9.3005
R7255 dvss.n2742 dvss.n2741 9.3005
R7256 dvss.n2740 dvss.n1740 9.3005
R7257 dvss.n1744 dvss.n1743 9.3005
R7258 dvss.n2734 dvss.n2733 9.3005
R7259 dvss.n2732 dvss.n2731 9.3005
R7260 dvss.n2730 dvss.n1747 9.3005
R7261 dvss.n2729 dvss.n2728 9.3005
R7262 dvss.n2727 dvss.n2726 9.3005
R7263 dvss.n2725 dvss.n1750 9.3005
R7264 dvss.n2724 dvss.n2723 9.3005
R7265 dvss.n2722 dvss.n2721 9.3005
R7266 dvss.n2720 dvss.n1753 9.3005
R7267 dvss.n2719 dvss.n2718 9.3005
R7268 dvss.n2717 dvss.n2716 9.3005
R7269 dvss.n1758 dvss.n1756 9.3005
R7270 dvss.n2711 dvss.n2710 9.3005
R7271 dvss.n2709 dvss.n2708 9.3005
R7272 dvss.n1764 dvss.n1761 9.3005
R7273 dvss.n2702 dvss.n2701 9.3005
R7274 dvss.n2700 dvss.n2699 9.3005
R7275 dvss.n1768 dvss.n1767 9.3005
R7276 dvss.n2694 dvss.n2693 9.3005
R7277 dvss.n2692 dvss.n2691 9.3005
R7278 dvss.n2690 dvss.n1771 9.3005
R7279 dvss.n1776 dvss.n1774 9.3005
R7280 dvss.n2684 dvss.n2683 9.3005
R7281 dvss.n1775 dvss.n168 9.3005
R7282 dvss.n3552 dvss.n3551 9.3005
R7283 dvss.n3553 dvss.n166 9.3005
R7284 dvss.n3568 dvss.n3567 9.3005
R7285 dvss.n3566 dvss.n167 9.3005
R7286 dvss.n3565 dvss.n3564 9.3005
R7287 dvss.n3563 dvss.n3562 9.3005
R7288 dvss.n3561 dvss.n3559 9.3005
R7289 dvss.n3560 dvss.n160 9.3005
R7290 dvss.n3577 dvss.n3576 9.3005
R7291 dvss.n3579 dvss.n157 9.3005
R7292 dvss.n3587 dvss.n3586 9.3005
R7293 dvss.n3585 dvss.n154 9.3005
R7294 dvss.n3594 dvss.n3593 9.3005
R7295 dvss.n3595 dvss.n149 9.3005
R7296 dvss.n3602 dvss.n3601 9.3005
R7297 dvss.n150 dvss.n144 9.3005
R7298 dvss.n3609 dvss.n3608 9.3005
R7299 dvss.n3610 dvss.n143 9.3005
R7300 dvss.n3620 dvss.n3619 9.3005
R7301 dvss.n3613 dvss.n139 9.3005
R7302 dvss.n3627 dvss.n3626 9.3005
R7303 dvss.n3628 dvss.n137 9.3005
R7304 dvss.n3633 dvss.n3632 9.3005
R7305 dvss.n3631 dvss.n138 9.3005
R7306 dvss.n3630 dvss.n133 9.3005
R7307 dvss.n3629 dvss.n131 9.3005
R7308 dvss.n3643 dvss.n3642 9.3005
R7309 dvss.n949 dvss.n861 9.3005
R7310 dvss.n956 dvss.n955 9.3005
R7311 dvss.n957 dvss.n763 9.3005
R7312 dvss.n963 dvss.n761 9.3005
R7313 dvss.n966 dvss.n965 9.3005
R7314 dvss.n972 dvss.n753 9.3005
R7315 dvss.n979 dvss.n978 9.3005
R7316 dvss.n755 dvss.n746 9.3005
R7317 dvss.n993 dvss.n992 9.3005
R7318 dvss.n984 dvss.n741 9.3005
R7319 dvss.n1001 dvss.n1000 9.3005
R7320 dvss.n738 dvss.n735 9.3005
R7321 dvss.n1017 dvss.n1016 9.3005
R7322 dvss.n1015 dvss.n726 9.3005
R7323 dvss.n1033 dvss.n1032 9.3005
R7324 dvss.n1031 dvss.n1030 9.3005
R7325 dvss.n1029 dvss.n718 9.3005
R7326 dvss.n1041 dvss.n1040 9.3005
R7327 dvss.n1042 dvss.n620 9.3005
R7328 dvss.n1043 dvss.n621 9.3005
R7329 dvss.n714 dvss.n622 9.3005
R7330 dvss.n1049 dvss.n1048 9.3005
R7331 dvss.n1052 dvss.n712 9.3005
R7332 dvss.n1059 dvss.n1058 9.3005
R7333 dvss.n1060 dvss.n631 9.3005
R7334 dvss.n1063 dvss.n632 9.3005
R7335 dvss.n1064 dvss.n633 9.3005
R7336 dvss.n1067 dvss.n1066 9.3005
R7337 dvss.n1065 dvss.n640 9.3005
R7338 dvss.n649 dvss.n641 9.3005
R7339 dvss.n1082 dvss.n642 9.3005
R7340 dvss.n1081 dvss.n1080 9.3005
R7341 dvss.n651 dvss.n650 9.3005
R7342 dvss.n707 dvss.n706 9.3005
R7343 dvss.n705 dvss.n704 9.3005
R7344 dvss.n703 dvss.n656 9.3005
R7345 dvss.n666 dvss.n664 9.3005
R7346 dvss.n693 dvss.n692 9.3005
R7347 dvss.n691 dvss.n690 9.3005
R7348 dvss.n1296 dvss.n565 9.3005
R7349 dvss.n1301 dvss.n1300 9.3005
R7350 dvss.n1302 dvss.n563 9.3005
R7351 dvss.n1318 dvss.n1317 9.3005
R7352 dvss.n1316 dvss.n1315 9.3005
R7353 dvss.n1314 dvss.n554 9.3005
R7354 dvss.n1328 dvss.n1327 9.3005
R7355 dvss.n1326 dvss.n552 9.3005
R7356 dvss.n1334 dvss.n548 9.3005
R7357 dvss.n1341 dvss.n1340 9.3005
R7358 dvss.n1347 dvss.n542 9.3005
R7359 dvss.n1354 dvss.n1353 9.3005
R7360 dvss.n1362 dvss.n538 9.3005
R7361 dvss.n1367 dvss.n1366 9.3005
R7362 dvss.n1365 dvss.n533 9.3005
R7363 dvss.n1378 dvss.n1377 9.3005
R7364 dvss.n1383 dvss.n529 9.3005
R7365 dvss.n1394 dvss.n1393 9.3005
R7366 dvss.n1392 dvss.n520 9.3005
R7367 dvss.n1410 dvss.n1409 9.3005
R7368 dvss.n1408 dvss.n1407 9.3005
R7369 dvss.n1406 dvss.n512 9.3005
R7370 dvss.n1417 dvss.n1416 9.3005
R7371 dvss.n1577 dvss.n1576 9.3005
R7372 dvss.n1575 dvss.n1574 9.3005
R7373 dvss.n1573 dvss.n1419 9.3005
R7374 dvss.n1572 dvss.n1571 9.3005
R7375 dvss.n1570 dvss.n1569 9.3005
R7376 dvss.n1568 dvss.n1424 9.3005
R7377 dvss.n1431 dvss.n1429 9.3005
R7378 dvss.n1564 dvss.n1563 9.3005
R7379 dvss.n1562 dvss.n1561 9.3005
R7380 dvss.n1499 dvss.n1434 9.3005
R7381 dvss.n1500 dvss.n1442 9.3005
R7382 dvss.n1555 dvss.n1554 9.3005
R7383 dvss.n1553 dvss.n1552 9.3005
R7384 dvss.n1551 dvss.n1445 9.3005
R7385 dvss.n1451 dvss.n1448 9.3005
R7386 dvss.n1544 dvss.n1543 9.3005
R7387 dvss.n1542 dvss.n1541 9.3005
R7388 dvss.n1540 dvss.n1454 9.3005
R7389 dvss.n1464 dvss.n1462 9.3005
R7390 dvss.n1530 dvss.n1529 9.3005
R7391 dvss.n1528 dvss.n1527 9.3005
R7392 dvss.n2886 dvss.n455 9.3005
R7393 dvss.n2891 dvss.n2890 9.3005
R7394 dvss.n2911 dvss.n2910 9.3005
R7395 dvss.n2909 dvss.n2908 9.3005
R7396 dvss.n2907 dvss.n2898 9.3005
R7397 dvss.n2906 dvss.n445 9.3005
R7398 dvss.n2920 dvss.n2919 9.3005
R7399 dvss.n2918 dvss.n443 9.3005
R7400 dvss.n2926 dvss.n439 9.3005
R7401 dvss.n2933 dvss.n2932 9.3005
R7402 dvss.n2939 dvss.n433 9.3005
R7403 dvss.n2946 dvss.n2945 9.3005
R7404 dvss.n2954 dvss.n429 9.3005
R7405 dvss.n2959 dvss.n2958 9.3005
R7406 dvss.n2957 dvss.n424 9.3005
R7407 dvss.n2970 dvss.n2969 9.3005
R7408 dvss.n2975 dvss.n420 9.3005
R7409 dvss.n2986 dvss.n2985 9.3005
R7410 dvss.n2984 dvss.n411 9.3005
R7411 dvss.n3003 dvss.n3002 9.3005
R7412 dvss.n3001 dvss.n3000 9.3005
R7413 dvss.n2999 dvss.n403 9.3005
R7414 dvss.n3010 dvss.n3009 9.3005
R7415 dvss.n3012 dvss.n3011 9.3005
R7416 dvss.n402 dvss.n396 9.3005
R7417 dvss.n3031 dvss.n3030 9.3005
R7418 dvss.n3029 dvss.n3028 9.3005
R7419 dvss.n3027 dvss.n3026 9.3005
R7420 dvss.n3039 dvss.n386 9.3005
R7421 dvss.n3046 dvss.n3045 9.3005
R7422 dvss.n3048 dvss.n3047 9.3005
R7423 dvss.n384 dvss.n381 9.3005
R7424 dvss.n3059 dvss.n374 9.3005
R7425 dvss.n3072 dvss.n3071 9.3005
R7426 dvss.n3074 dvss.n3073 9.3005
R7427 dvss.n3065 dvss.n364 9.3005
R7428 dvss.n3084 dvss.n3083 9.3005
R7429 dvss.n3086 dvss.n3085 9.3005
R7430 dvss.n3091 dvss.n358 9.3005
R7431 dvss.n3098 dvss.n3097 9.3005
R7432 dvss.n3105 dvss.n348 9.3005
R7433 dvss.n3120 dvss.n3119 9.3005
R7434 dvss.n3118 dvss.n3117 9.3005
R7435 dvss.n3116 dvss.n351 9.3005
R7436 dvss.n3126 dvss.n338 9.3005
R7437 dvss.n3131 dvss.n3130 9.3005
R7438 dvss.n3129 dvss.n326 9.3005
R7439 dvss.n3145 dvss.n3144 9.3005
R7440 dvss.n3143 dvss.n327 9.3005
R7441 dvss.n3142 dvss.n321 9.3005
R7442 dvss.n3153 dvss.n3152 9.3005
R7443 dvss.n3151 dvss.n319 9.3005
R7444 dvss.n3165 dvss.n316 9.3005
R7445 dvss.n3160 dvss.n311 9.3005
R7446 dvss.n3177 dvss.n3176 9.3005
R7447 dvss.n3179 dvss.n3178 9.3005
R7448 dvss.n3187 dvss.n306 9.3005
R7449 dvss.n309 dvss.n300 9.3005
R7450 dvss.n3200 dvss.n3199 9.3005
R7451 dvss.n3202 dvss.n3201 9.3005
R7452 dvss.n3207 dvss.n294 9.3005
R7453 dvss.n3214 dvss.n3213 9.3005
R7454 dvss.n3221 dvss.n284 9.3005
R7455 dvss.n3236 dvss.n3235 9.3005
R7456 dvss.n3234 dvss.n3233 9.3005
R7457 dvss.n3232 dvss.n287 9.3005
R7458 dvss.n3242 dvss.n274 9.3005
R7459 dvss.n3247 dvss.n3246 9.3005
R7460 dvss.n3245 dvss.n262 9.3005
R7461 dvss.n3261 dvss.n3260 9.3005
R7462 dvss.n3259 dvss.n263 9.3005
R7463 dvss.n3258 dvss.n257 9.3005
R7464 dvss.n3268 dvss.n3267 9.3005
R7465 dvss.n3274 dvss.n254 9.3005
R7466 dvss.n3284 dvss.n3283 9.3005
R7467 dvss.n3278 dvss.n247 9.3005
R7468 dvss.n3293 dvss.n3292 9.3005
R7469 dvss.n3294 dvss.n243 9.3005
R7470 dvss.n3306 dvss.n3305 9.3005
R7471 dvss.n3304 dvss.n3303 9.3005
R7472 dvss.n3302 dvss.n234 9.3005
R7473 dvss.n3318 dvss.n3317 9.3005
R7474 dvss.n3323 dvss.n230 9.3005
R7475 dvss.n3334 dvss.n3333 9.3005
R7476 dvss.n3332 dvss.n221 9.3005
R7477 dvss.n3350 dvss.n3349 9.3005
R7478 dvss.n3348 dvss.n3347 9.3005
R7479 dvss.n3346 dvss.n213 9.3005
R7480 dvss.n3357 dvss.n3356 9.3005
R7481 dvss.n3543 dvss.n3542 9.3005
R7482 dvss.n3541 dvss.n3540 9.3005
R7483 dvss.n3539 dvss.n3359 9.3005
R7484 dvss.n3538 dvss.n3537 9.3005
R7485 dvss.n3536 dvss.n3535 9.3005
R7486 dvss.n3534 dvss.n3364 9.3005
R7487 dvss.n3371 dvss.n3369 9.3005
R7488 dvss.n3530 dvss.n3529 9.3005
R7489 dvss.n3528 dvss.n3527 9.3005
R7490 dvss.n3426 dvss.n3374 9.3005
R7491 dvss.n3427 dvss.n3382 9.3005
R7492 dvss.n3521 dvss.n3520 9.3005
R7493 dvss.n3519 dvss.n3518 9.3005
R7494 dvss.n3517 dvss.n3385 9.3005
R7495 dvss.n3391 dvss.n3388 9.3005
R7496 dvss.n3510 dvss.n3509 9.3005
R7497 dvss.n3508 dvss.n3507 9.3005
R7498 dvss.n3506 dvss.n3394 9.3005
R7499 dvss.n3473 dvss.n3399 9.3005
R7500 dvss.n3475 dvss.n3474 9.3005
R7501 dvss.n3418 dvss.n3413 9.3005
R7502 dvss.n3417 dvss.n3406 9.3005
R7503 dvss.n3494 dvss.n3493 9.3005
R7504 dvss.n3492 dvss.n3491 9.3005
R7505 dvss.n3490 dvss.n124 9.3005
R7506 dvss.n3647 dvss.n3646 9.3005
R7507 dvss.n2663 dvss.n1966 9.3005
R7508 dvss.n2662 dvss.n2661 9.3005
R7509 dvss.n2660 dvss.n2659 9.3005
R7510 dvss.n2645 dvss.n2644 9.3005
R7511 dvss.n2646 dvss.n2645 9.3005
R7512 dvss.n2637 dvss.n2636 9.3005
R7513 dvss.n2638 dvss.n2637 9.3005
R7514 dvss.n2626 dvss.n2625 9.3005
R7515 dvss.n2627 dvss.n2626 9.3005
R7516 dvss.n2592 dvss.n2591 9.3005
R7517 dvss.n2593 dvss.n2592 9.3005
R7518 dvss.n2601 dvss.n2599 9.3005
R7519 dvss.n2602 dvss.n2601 9.3005
R7520 dvss.n2609 dvss.n2607 9.3005
R7521 dvss.n2610 dvss.n2609 9.3005
R7522 dvss.n2579 dvss.n2578 9.3005
R7523 dvss.n2580 dvss.n2579 9.3005
R7524 dvss.n2545 dvss.n2544 9.3005
R7525 dvss.n2546 dvss.n2545 9.3005
R7526 dvss.n2554 dvss.n2552 9.3005
R7527 dvss.n2555 dvss.n2554 9.3005
R7528 dvss.n2562 dvss.n2560 9.3005
R7529 dvss.n2563 dvss.n2562 9.3005
R7530 dvss.n2532 dvss.n2531 9.3005
R7531 dvss.n2533 dvss.n2532 9.3005
R7532 dvss.n2498 dvss.n2497 9.3005
R7533 dvss.n2499 dvss.n2498 9.3005
R7534 dvss.n2507 dvss.n2505 9.3005
R7535 dvss.n2508 dvss.n2507 9.3005
R7536 dvss.n2515 dvss.n2513 9.3005
R7537 dvss.n2516 dvss.n2515 9.3005
R7538 dvss.n2485 dvss.n2484 9.3005
R7539 dvss.n2486 dvss.n2485 9.3005
R7540 dvss.n2451 dvss.n2450 9.3005
R7541 dvss.n2452 dvss.n2451 9.3005
R7542 dvss.n2460 dvss.n2458 9.3005
R7543 dvss.n2461 dvss.n2460 9.3005
R7544 dvss.n2468 dvss.n2466 9.3005
R7545 dvss.n2469 dvss.n2468 9.3005
R7546 dvss.n2438 dvss.n2437 9.3005
R7547 dvss.n2439 dvss.n2438 9.3005
R7548 dvss.n2404 dvss.n2403 9.3005
R7549 dvss.n2405 dvss.n2404 9.3005
R7550 dvss.n2413 dvss.n2411 9.3005
R7551 dvss.n2414 dvss.n2413 9.3005
R7552 dvss.n2421 dvss.n2419 9.3005
R7553 dvss.n2422 dvss.n2421 9.3005
R7554 dvss.n2391 dvss.n2390 9.3005
R7555 dvss.n2392 dvss.n2391 9.3005
R7556 dvss.n2357 dvss.n2356 9.3005
R7557 dvss.n2358 dvss.n2357 9.3005
R7558 dvss.n2366 dvss.n2364 9.3005
R7559 dvss.n2367 dvss.n2366 9.3005
R7560 dvss.n2374 dvss.n2372 9.3005
R7561 dvss.n2375 dvss.n2374 9.3005
R7562 dvss.n2344 dvss.n2343 9.3005
R7563 dvss.n2345 dvss.n2344 9.3005
R7564 dvss.n2310 dvss.n2309 9.3005
R7565 dvss.n2311 dvss.n2310 9.3005
R7566 dvss.n2319 dvss.n2317 9.3005
R7567 dvss.n2320 dvss.n2319 9.3005
R7568 dvss.n2327 dvss.n2325 9.3005
R7569 dvss.n2328 dvss.n2327 9.3005
R7570 dvss.n2297 dvss.n2296 9.3005
R7571 dvss.n2298 dvss.n2297 9.3005
R7572 dvss.n3708 dvss.n3707 9.3005
R7573 dvss.n3709 dvss.n3708 9.3005
R7574 dvss.n3717 dvss.n3715 9.3005
R7575 dvss.n3718 dvss.n3717 9.3005
R7576 dvss.n3725 dvss.n3723 9.3005
R7577 dvss.n3726 dvss.n3725 9.3005
R7578 dvss.n3695 dvss.n3694 9.3005
R7579 dvss.n3696 dvss.n3695 9.3005
R7580 dvss.n3661 dvss.n3660 9.3005
R7581 dvss.n3662 dvss.n3661 9.3005
R7582 dvss.n3670 dvss.n3668 9.3005
R7583 dvss.n3671 dvss.n3670 9.3005
R7584 dvss.n3678 dvss.n3676 9.3005
R7585 dvss.n3679 dvss.n3678 9.3005
R7586 dvss.n2657 dvss.n1969 9.3005
R7587 dvss.n2656 dvss.n2655 9.3005
R7588 dvss.n2654 dvss.n2653 9.3005
R7589 dvss.n2652 dvss.n1974 9.3005
R7590 dvss.n2651 dvss.n2650 9.3005
R7591 dvss.n2649 dvss.n2648 9.3005
R7592 dvss.n2647 dvss.n1977 9.3005
R7593 dvss.n2643 dvss.n2642 9.3005
R7594 dvss.n2641 dvss.n2640 9.3005
R7595 dvss.n2639 dvss.n1985 9.3005
R7596 dvss.n1990 dvss.n1989 9.3005
R7597 dvss.n2635 dvss.n2634 9.3005
R7598 dvss.n2633 dvss.n2632 9.3005
R7599 dvss.n2631 dvss.n2630 9.3005
R7600 dvss.n2629 dvss.n2628 9.3005
R7601 dvss.n2000 dvss.n1997 9.3005
R7602 dvss.n2624 dvss.n2623 9.3005
R7603 dvss.n2622 dvss.n2621 9.3005
R7604 dvss.n2620 dvss.n2003 9.3005
R7605 dvss.n2619 dvss.n2618 9.3005
R7606 dvss.n2617 dvss.n2616 9.3005
R7607 dvss.n2615 dvss.n2008 9.3005
R7608 dvss.n2614 dvss.n2613 9.3005
R7609 dvss.n2612 dvss.n2611 9.3005
R7610 dvss.n2013 dvss.n2011 9.3005
R7611 dvss.n2606 dvss.n2605 9.3005
R7612 dvss.n2604 dvss.n2603 9.3005
R7613 dvss.n2019 dvss.n2018 9.3005
R7614 dvss.n2598 dvss.n2597 9.3005
R7615 dvss.n2596 dvss.n2595 9.3005
R7616 dvss.n2594 dvss.n2022 9.3005
R7617 dvss.n2590 dvss.n2589 9.3005
R7618 dvss.n2588 dvss.n2587 9.3005
R7619 dvss.n2586 dvss.n2027 9.3005
R7620 dvss.n2585 dvss.n2584 9.3005
R7621 dvss.n2583 dvss.n2582 9.3005
R7622 dvss.n2581 dvss.n2030 9.3005
R7623 dvss.n2036 dvss.n2033 9.3005
R7624 dvss.n2577 dvss.n2576 9.3005
R7625 dvss.n2575 dvss.n2574 9.3005
R7626 dvss.n2573 dvss.n2039 9.3005
R7627 dvss.n2572 dvss.n2571 9.3005
R7628 dvss.n2570 dvss.n2569 9.3005
R7629 dvss.n2568 dvss.n2044 9.3005
R7630 dvss.n2567 dvss.n2566 9.3005
R7631 dvss.n2565 dvss.n2564 9.3005
R7632 dvss.n2049 dvss.n2047 9.3005
R7633 dvss.n2559 dvss.n2558 9.3005
R7634 dvss.n2557 dvss.n2556 9.3005
R7635 dvss.n2055 dvss.n2054 9.3005
R7636 dvss.n2551 dvss.n2550 9.3005
R7637 dvss.n2549 dvss.n2548 9.3005
R7638 dvss.n2547 dvss.n2058 9.3005
R7639 dvss.n2543 dvss.n2542 9.3005
R7640 dvss.n2541 dvss.n2540 9.3005
R7641 dvss.n2539 dvss.n2063 9.3005
R7642 dvss.n2538 dvss.n2537 9.3005
R7643 dvss.n2536 dvss.n2535 9.3005
R7644 dvss.n2534 dvss.n2066 9.3005
R7645 dvss.n2072 dvss.n2069 9.3005
R7646 dvss.n2530 dvss.n2529 9.3005
R7647 dvss.n2528 dvss.n2527 9.3005
R7648 dvss.n2526 dvss.n2075 9.3005
R7649 dvss.n2525 dvss.n2524 9.3005
R7650 dvss.n2523 dvss.n2522 9.3005
R7651 dvss.n2521 dvss.n2080 9.3005
R7652 dvss.n2520 dvss.n2519 9.3005
R7653 dvss.n2518 dvss.n2517 9.3005
R7654 dvss.n2085 dvss.n2083 9.3005
R7655 dvss.n2512 dvss.n2511 9.3005
R7656 dvss.n2510 dvss.n2509 9.3005
R7657 dvss.n2091 dvss.n2090 9.3005
R7658 dvss.n2504 dvss.n2503 9.3005
R7659 dvss.n2502 dvss.n2501 9.3005
R7660 dvss.n2500 dvss.n2094 9.3005
R7661 dvss.n2496 dvss.n2495 9.3005
R7662 dvss.n2494 dvss.n2493 9.3005
R7663 dvss.n2492 dvss.n2099 9.3005
R7664 dvss.n2491 dvss.n2490 9.3005
R7665 dvss.n2489 dvss.n2488 9.3005
R7666 dvss.n2487 dvss.n2102 9.3005
R7667 dvss.n2108 dvss.n2105 9.3005
R7668 dvss.n2483 dvss.n2482 9.3005
R7669 dvss.n2481 dvss.n2480 9.3005
R7670 dvss.n2479 dvss.n2111 9.3005
R7671 dvss.n2478 dvss.n2477 9.3005
R7672 dvss.n2476 dvss.n2475 9.3005
R7673 dvss.n2474 dvss.n2116 9.3005
R7674 dvss.n2473 dvss.n2472 9.3005
R7675 dvss.n2471 dvss.n2470 9.3005
R7676 dvss.n2121 dvss.n2119 9.3005
R7677 dvss.n2465 dvss.n2464 9.3005
R7678 dvss.n2463 dvss.n2462 9.3005
R7679 dvss.n2127 dvss.n2126 9.3005
R7680 dvss.n2457 dvss.n2456 9.3005
R7681 dvss.n2455 dvss.n2454 9.3005
R7682 dvss.n2453 dvss.n2130 9.3005
R7683 dvss.n2449 dvss.n2448 9.3005
R7684 dvss.n2447 dvss.n2446 9.3005
R7685 dvss.n2445 dvss.n2135 9.3005
R7686 dvss.n2444 dvss.n2443 9.3005
R7687 dvss.n2442 dvss.n2441 9.3005
R7688 dvss.n2440 dvss.n2138 9.3005
R7689 dvss.n2144 dvss.n2141 9.3005
R7690 dvss.n2436 dvss.n2435 9.3005
R7691 dvss.n2434 dvss.n2433 9.3005
R7692 dvss.n2432 dvss.n2147 9.3005
R7693 dvss.n2431 dvss.n2430 9.3005
R7694 dvss.n2429 dvss.n2428 9.3005
R7695 dvss.n2427 dvss.n2152 9.3005
R7696 dvss.n2426 dvss.n2425 9.3005
R7697 dvss.n2424 dvss.n2423 9.3005
R7698 dvss.n2157 dvss.n2155 9.3005
R7699 dvss.n2418 dvss.n2417 9.3005
R7700 dvss.n2416 dvss.n2415 9.3005
R7701 dvss.n2163 dvss.n2162 9.3005
R7702 dvss.n2410 dvss.n2409 9.3005
R7703 dvss.n2408 dvss.n2407 9.3005
R7704 dvss.n2406 dvss.n2166 9.3005
R7705 dvss.n2402 dvss.n2401 9.3005
R7706 dvss.n2400 dvss.n2399 9.3005
R7707 dvss.n2398 dvss.n2171 9.3005
R7708 dvss.n2397 dvss.n2396 9.3005
R7709 dvss.n2395 dvss.n2394 9.3005
R7710 dvss.n2393 dvss.n2174 9.3005
R7711 dvss.n2180 dvss.n2177 9.3005
R7712 dvss.n2389 dvss.n2388 9.3005
R7713 dvss.n2387 dvss.n2386 9.3005
R7714 dvss.n2385 dvss.n2183 9.3005
R7715 dvss.n2384 dvss.n2383 9.3005
R7716 dvss.n2382 dvss.n2381 9.3005
R7717 dvss.n2380 dvss.n2188 9.3005
R7718 dvss.n2379 dvss.n2378 9.3005
R7719 dvss.n2377 dvss.n2376 9.3005
R7720 dvss.n2194 dvss.n2192 9.3005
R7721 dvss.n2371 dvss.n2370 9.3005
R7722 dvss.n2369 dvss.n2368 9.3005
R7723 dvss.n2197 dvss.n2196 9.3005
R7724 dvss.n2363 dvss.n2362 9.3005
R7725 dvss.n2361 dvss.n2360 9.3005
R7726 dvss.n2359 dvss.n2200 9.3005
R7727 dvss.n2355 dvss.n2354 9.3005
R7728 dvss.n2353 dvss.n2352 9.3005
R7729 dvss.n2351 dvss.n2203 9.3005
R7730 dvss.n2350 dvss.n2349 9.3005
R7731 dvss.n2348 dvss.n2347 9.3005
R7732 dvss.n2346 dvss.n2206 9.3005
R7733 dvss.n2210 dvss.n2209 9.3005
R7734 dvss.n2342 dvss.n2341 9.3005
R7735 dvss.n2340 dvss.n2339 9.3005
R7736 dvss.n2338 dvss.n2213 9.3005
R7737 dvss.n2337 dvss.n2336 9.3005
R7738 dvss.n2335 dvss.n2334 9.3005
R7739 dvss.n2333 dvss.n2216 9.3005
R7740 dvss.n2332 dvss.n2331 9.3005
R7741 dvss.n2330 dvss.n2329 9.3005
R7742 dvss.n2248 dvss.n2246 9.3005
R7743 dvss.n2324 dvss.n2323 9.3005
R7744 dvss.n2322 dvss.n2321 9.3005
R7745 dvss.n2252 dvss.n2251 9.3005
R7746 dvss.n2316 dvss.n2315 9.3005
R7747 dvss.n2314 dvss.n2313 9.3005
R7748 dvss.n2312 dvss.n2255 9.3005
R7749 dvss.n2308 dvss.n2307 9.3005
R7750 dvss.n2306 dvss.n2305 9.3005
R7751 dvss.n2304 dvss.n2258 9.3005
R7752 dvss.n2303 dvss.n2302 9.3005
R7753 dvss.n2301 dvss.n2300 9.3005
R7754 dvss.n2299 dvss.n2292 9.3005
R7755 dvss.n2295 dvss.n68 9.3005
R7756 dvss.n3740 dvss.n3739 9.3005
R7757 dvss.n3738 dvss.n3737 9.3005
R7758 dvss.n3736 dvss.n71 9.3005
R7759 dvss.n3735 dvss.n3734 9.3005
R7760 dvss.n3733 dvss.n3732 9.3005
R7761 dvss.n3731 dvss.n74 9.3005
R7762 dvss.n3730 dvss.n3729 9.3005
R7763 dvss.n3728 dvss.n3727 9.3005
R7764 dvss.n79 dvss.n77 9.3005
R7765 dvss.n3722 dvss.n3721 9.3005
R7766 dvss.n3720 dvss.n3719 9.3005
R7767 dvss.n83 dvss.n82 9.3005
R7768 dvss.n3714 dvss.n3713 9.3005
R7769 dvss.n3712 dvss.n3711 9.3005
R7770 dvss.n3710 dvss.n86 9.3005
R7771 dvss.n3706 dvss.n3705 9.3005
R7772 dvss.n3704 dvss.n3703 9.3005
R7773 dvss.n3702 dvss.n89 9.3005
R7774 dvss.n3701 dvss.n3700 9.3005
R7775 dvss.n3699 dvss.n3698 9.3005
R7776 dvss.n3697 dvss.n92 9.3005
R7777 dvss.n96 dvss.n95 9.3005
R7778 dvss.n3693 dvss.n3692 9.3005
R7779 dvss.n3691 dvss.n3690 9.3005
R7780 dvss.n3689 dvss.n99 9.3005
R7781 dvss.n3688 dvss.n3687 9.3005
R7782 dvss.n3686 dvss.n3685 9.3005
R7783 dvss.n3684 dvss.n102 9.3005
R7784 dvss.n3683 dvss.n3682 9.3005
R7785 dvss.n3681 dvss.n3680 9.3005
R7786 dvss.n107 dvss.n105 9.3005
R7787 dvss.n3675 dvss.n3674 9.3005
R7788 dvss.n3673 dvss.n3672 9.3005
R7789 dvss.n111 dvss.n110 9.3005
R7790 dvss.n3667 dvss.n3666 9.3005
R7791 dvss.n3665 dvss.n3664 9.3005
R7792 dvss.n3663 dvss.n114 9.3005
R7793 dvss.n3659 dvss.n3658 9.3005
R7794 dvss.n3657 dvss.n3656 9.3005
R7795 dvss.n3655 dvss.n117 9.3005
R7796 dvss.n3654 dvss.n3653 9.3005
R7797 dvss.n3745 dvss.n3 9.3005
R7798 dvss.n3747 dvss.n3746 9.3005
R7799 dvss.n3748 dvss.n0 9.3005
R7800 dvss.n3751 dvss.n3750 9.3005
R7801 dvss.n47 dvss.n1 9.3005
R7802 dvss.n27 dvss.n26 9.3005
R7803 dvss.n29 dvss.n21 9.3005
R7804 dvss.n33 dvss.n32 9.3005
R7805 dvss.n34 dvss.n20 9.3005
R7806 dvss.n36 dvss.n35 9.3005
R7807 dvss.n38 dvss.n18 9.3005
R7808 dvss.n42 dvss.n41 9.3005
R7809 dvss.n43 dvss.n15 9.3005
R7810 dvss.n55 dvss.n54 9.3005
R7811 dvss.n53 dvss.n52 9.3005
R7812 dvss.n50 dvss.n44 9.3005
R7813 dvss.n49 dvss.n48 9.3005
R7814 dvss.n943 dvss.t316 9.09947
R7815 dvss.n1988 dvss.n1986 8.56999
R7816 dvss.n3695 dvss.n94 8.54791
R7817 dvss.n2297 dvss.n2294 8.54791
R7818 dvss.n2344 dvss.n2208 8.54791
R7819 dvss.n2391 dvss.n2176 8.54791
R7820 dvss.n2438 dvss.n2140 8.54791
R7821 dvss.n2485 dvss.n2104 8.54791
R7822 dvss.n2532 dvss.n2068 8.54791
R7823 dvss.n2579 dvss.n2032 8.54791
R7824 dvss.n2626 dvss.n1999 8.54791
R7825 dvss.n3532 dvss.n3368 8.54791
R7826 dvss.n3272 dvss.n3271 8.54791
R7827 dvss.n3157 dvss.n3156 8.54791
R7828 dvss.n3043 dvss.n3042 8.54791
R7829 dvss.n2924 dvss.n2923 8.54791
R7830 dvss.n1566 dvss.n1428 8.54791
R7831 dvss.n1332 dvss.n1331 8.54791
R7832 dvss.n1056 dvss.n1054 8.54791
R7833 dvss.n953 dvss.n951 8.54791
R7834 dvss.n1978 dvss 8.48432
R7835 dvss.n94 dvss 8.43944
R7836 dvss.n2294 dvss 8.43944
R7837 dvss.n2208 dvss 8.43944
R7838 dvss.n2176 dvss 8.43944
R7839 dvss.n2140 dvss 8.43944
R7840 dvss.n2104 dvss 8.43944
R7841 dvss.n2068 dvss 8.43944
R7842 dvss.n2032 dvss 8.43944
R7843 dvss.n1999 dvss 8.43944
R7844 dvss.n3368 dvss 8.43944
R7845 dvss.n3271 dvss 8.43944
R7846 dvss.n3156 dvss 8.43944
R7847 dvss.n3042 dvss 8.43944
R7848 dvss.n2923 dvss 8.43944
R7849 dvss.n1428 dvss 8.43944
R7850 dvss.n1331 dvss 8.43944
R7851 dvss.n1054 dvss 8.43944
R7852 dvss.n951 dvss 8.43944
R7853 dvss.n38 dvss.n37 8.2416
R7854 dvss.n901 dvss.t78 8.21389
R7855 dvss.n37 dvss.n36 7.89091
R7856 dvss.n904 dvss.t475 7.79961
R7857 dvss.n2637 dvss.n1988 7.37677
R7858 dvss.n3397 dvss 6.4005
R7859 dvss.n3327 dvss 6.4005
R7860 dvss.n3216 dvss 6.4005
R7861 dvss.n3100 dvss 6.4005
R7862 dvss.n2979 dvss 6.4005
R7863 dvss.n1460 dvss 6.4005
R7864 dvss.n1387 dvss 6.4005
R7865 dvss.n662 dvss 6.4005
R7866 dvss.n1010 dvss 6.4005
R7867 dvss.n3611 dvss 6.4005
R7868 dvss.n1772 dvss 6.4005
R7869 dvss.n1741 dvss 6.4005
R7870 dvss.n1710 dvss 6.4005
R7871 dvss.n1679 dvss 6.4005
R7872 dvss.n474 dvss 6.4005
R7873 dvss.n1206 dvss 6.4005
R7874 dvss.n584 dvss 6.4005
R7875 dvss.n816 dvss 6.4005
R7876 dvss.n25 dvss.n24 5.87299
R7877 dvss.n767 dvss 5.69343
R7878 dvss.n3504 dvss 5.45235
R7879 dvss.n3330 dvss 5.45235
R7880 dvss.n3219 dvss 5.45235
R7881 dvss.n3103 dvss 5.45235
R7882 dvss.n2982 dvss 5.45235
R7883 dvss.n1538 dvss 5.45235
R7884 dvss.n1390 dvss 5.45235
R7885 dvss.n701 dvss 5.45235
R7886 dvss.n1013 dvss 5.45235
R7887 dvss.n3617 dvss 5.45235
R7888 dvss.n2688 dvss 5.45235
R7889 dvss.n2738 dvss 5.45235
R7890 dvss.n2788 dvss 5.45235
R7891 dvss.n2838 dvss 5.45235
R7892 dvss.n1644 dvss 5.45235
R7893 dvss.n1248 dvss 5.45235
R7894 dvss.n1171 dvss 5.45235
R7895 dvss.n815 dvss 5.45235
R7896 dvss.n31 dvss.n20 5.43612
R7897 dvss.n41 dvss.n40 5.08543
R7898 dvss dvss.n3742 4.88201
R7899 dvss.n941 dvss.t255 3.90006
R7900 dvss dvss.n3741 3.78956
R7901 dvss.n3670 dvss.n106 3.68864
R7902 dvss.n3717 dvss.n78 3.68864
R7903 dvss.n2319 dvss.n2247 3.68864
R7904 dvss.n2366 dvss.n2193 3.68864
R7905 dvss.n2413 dvss.n2156 3.68864
R7906 dvss.n2460 dvss.n2120 3.68864
R7907 dvss.n2507 dvss.n2084 3.68864
R7908 dvss.n2554 dvss.n2048 3.68864
R7909 dvss.n2601 dvss.n2012 3.68864
R7910 dvss.n3500 dvss.n3497 3.68864
R7911 dvss.n3353 dvss.n3352 3.68864
R7912 dvss.n3239 dvss.n3238 3.68864
R7913 dvss.n3123 dvss.n3122 3.68864
R7914 dvss.n3006 dvss.n3005 3.68864
R7915 dvss.n1534 dvss.n457 3.68864
R7916 dvss.n1413 dvss.n1412 3.68864
R7917 dvss.n697 dvss.n567 3.68864
R7918 dvss.n1036 dvss.n1035 3.68864
R7919 dvss.n3742 dvss.n67 3.60119
R7920 dvss.n767 dvss 3.53935
R7921 dvss.n1986 dvss 3.25474
R7922 dvss.n3645 dvss 2.94111
R7923 dvss.n3504 dvss.n3503 2.84494
R7924 dvss.n3330 dvss.n3329 2.84494
R7925 dvss.n3219 dvss.n3218 2.84494
R7926 dvss.n3103 dvss.n3102 2.84494
R7927 dvss.n2982 dvss.n2981 2.84494
R7928 dvss.n1538 dvss.n1537 2.84494
R7929 dvss.n1390 dvss.n1389 2.84494
R7930 dvss.n701 dvss.n700 2.84494
R7931 dvss.n1013 dvss.n1012 2.84494
R7932 dvss.n3617 dvss.n3616 2.84494
R7933 dvss.n2688 dvss.n2687 2.84494
R7934 dvss.n2738 dvss.n2737 2.84494
R7935 dvss.n2788 dvss.n2787 2.84494
R7936 dvss.n2838 dvss.n2837 2.84494
R7937 dvss.n1645 dvss.n1644 2.84494
R7938 dvss.n1248 dvss.n1247 2.84494
R7939 dvss.n1172 dvss.n1171 2.84494
R7940 dvss.n815 dvss.n814 2.84494
R7941 dvss.n29 dvss.n28 2.63064
R7942 dvss.n3503 dvss 2.60791
R7943 dvss.n3329 dvss 2.60791
R7944 dvss.n3218 dvss 2.60791
R7945 dvss.n3102 dvss 2.60791
R7946 dvss.n2981 dvss 2.60791
R7947 dvss.n1537 dvss 2.60791
R7948 dvss.n1389 dvss 2.60791
R7949 dvss.n700 dvss 2.60791
R7950 dvss.n1012 dvss 2.60791
R7951 dvss.n3616 dvss 2.60791
R7952 dvss.n2687 dvss 2.60791
R7953 dvss.n2737 dvss 2.60791
R7954 dvss.n2787 dvss 2.60791
R7955 dvss.n2837 dvss 2.60791
R7956 dvss.n1645 dvss 2.60791
R7957 dvss.n1247 dvss 2.60791
R7958 dvss.n1172 dvss 2.60791
R7959 dvss.n814 dvss 2.60791
R7960 dvss.t308 dvss.t78 2.57737
R7961 dvss.n916 dvss 2.49542
R7962 dvss.n911 dvss 2.49542
R7963 dvss.n55 dvss.n17 2.27995
R7964 dvss.n46 dvss.n1 2.27995
R7965 dvss.n8 dvss.n7 2.17238
R7966 dvss.n885 dvss 2.16773
R7967 dvss.n2658 dvss 2.16773
R7968 dvss.n3515 dvss 1.84457
R7969 dvss dvss.n3514 1.84457
R7970 dvss.n3514 dvss 1.84457
R7971 dvss.n3320 dvss 1.84457
R7972 dvss.n3299 dvss 1.84457
R7973 dvss.n3299 dvss 1.84457
R7974 dvss.n3204 dvss 1.84457
R7975 dvss.n3184 dvss 1.84457
R7976 dvss.n3184 dvss 1.84457
R7977 dvss.n3088 dvss 1.84457
R7978 dvss.n3064 dvss 1.84457
R7979 dvss.n3064 dvss 1.84457
R7980 dvss.n2972 dvss 1.84457
R7981 dvss.n2951 dvss 1.84457
R7982 dvss.n2951 dvss 1.84457
R7983 dvss.n1549 dvss 1.84457
R7984 dvss dvss.n1548 1.84457
R7985 dvss.n1548 dvss 1.84457
R7986 dvss.n1380 dvss 1.84457
R7987 dvss.n1359 dvss 1.84457
R7988 dvss.n1359 dvss 1.84457
R7989 dvss.n1078 dvss 1.84457
R7990 dvss dvss.n1077 1.84457
R7991 dvss.n1077 dvss 1.84457
R7992 dvss.n997 dvss 1.84457
R7993 dvss dvss.n996 1.84457
R7994 dvss.n996 dvss 1.84457
R7995 dvss.n3599 dvss 1.84457
R7996 dvss dvss.n3598 1.84457
R7997 dvss.n3598 dvss 1.84457
R7998 dvss.n2697 dvss 1.84457
R7999 dvss dvss.n2696 1.84457
R8000 dvss.n2696 dvss 1.84457
R8001 dvss.n2747 dvss 1.84457
R8002 dvss dvss.n2746 1.84457
R8003 dvss.n2746 dvss 1.84457
R8004 dvss.n2797 dvss 1.84457
R8005 dvss dvss.n2796 1.84457
R8006 dvss.n2796 dvss 1.84457
R8007 dvss.n2847 dvss 1.84457
R8008 dvss dvss.n2846 1.84457
R8009 dvss.n2846 dvss 1.84457
R8010 dvss.n1630 dvss 1.84457
R8011 dvss dvss.n1629 1.84457
R8012 dvss.n1629 dvss 1.84457
R8013 dvss.n1257 dvss 1.84457
R8014 dvss dvss.n1256 1.84457
R8015 dvss.n1256 dvss 1.84457
R8016 dvss.n1157 dvss 1.84457
R8017 dvss dvss.n1156 1.84457
R8018 dvss.n1156 dvss 1.84457
R8019 dvss.n801 dvss 1.84457
R8020 dvss dvss.n799 1.84457
R8021 dvss.n799 dvss 1.84457
R8022 dvss.n3645 dvss.n3644 1.5923
R8023 dvss.n56 dvss.n15 1.57858
R8024 dvss.n3750 dvss.n3749 1.40324
R8025 dvss.n3525 dvss.n3378 1.34003
R8026 dvss.n3523 dvss.n3380 1.34003
R8027 dvss.n3513 dvss.n3380 1.34003
R8028 dvss.n3281 dvss.n3280 1.34003
R8029 dvss.n3298 dvss.n3296 1.34003
R8030 dvss.n3300 dvss.n3298 1.34003
R8031 dvss.n3163 dvss.n3162 1.34003
R8032 dvss.n3183 dvss.n3181 1.34003
R8033 dvss.n3185 dvss.n3183 1.34003
R8034 dvss.n3061 dvss.n377 1.34003
R8035 dvss.n3069 dvss.n3068 1.34003
R8036 dvss.n3068 dvss.n3067 1.34003
R8037 dvss.n2937 dvss.n2936 1.34003
R8038 dvss.n2950 dvss.n2948 1.34003
R8039 dvss.n2952 dvss.n2950 1.34003
R8040 dvss.n1559 dvss.n1438 1.34003
R8041 dvss.n1557 dvss.n1440 1.34003
R8042 dvss.n1547 dvss.n1440 1.34003
R8043 dvss.n1345 dvss.n1344 1.34003
R8044 dvss.n1358 dvss.n1356 1.34003
R8045 dvss.n1360 dvss.n1358 1.34003
R8046 dvss.n1069 dvss.n711 1.34003
R8047 dvss.n1074 dvss.n1072 1.34003
R8048 dvss.n1076 dvss.n1074 1.34003
R8049 dvss.n974 dvss.n757 1.34003
R8050 dvss.n976 dvss.n744 1.34003
R8051 dvss.n995 dvss.n744 1.34003
R8052 dvss.n3581 dvss.n159 1.34003
R8053 dvss.n3583 dvss.n153 1.34003
R8054 dvss.n3597 dvss.n153 1.34003
R8055 dvss.n2714 dvss.n2713 1.34003
R8056 dvss.n2706 dvss.n2705 1.34003
R8057 dvss.n2705 dvss.n2704 1.34003
R8058 dvss.n2764 dvss.n2763 1.34003
R8059 dvss.n2756 dvss.n2755 1.34003
R8060 dvss.n2755 dvss.n2754 1.34003
R8061 dvss.n2814 dvss.n2813 1.34003
R8062 dvss.n2806 dvss.n2805 1.34003
R8063 dvss.n2805 dvss.n2804 1.34003
R8064 dvss.n2864 dvss.n2863 1.34003
R8065 dvss.n2856 dvss.n2855 1.34003
R8066 dvss.n2855 dvss.n2854 1.34003
R8067 dvss.n1613 dvss.n491 1.34003
R8068 dvss.n1615 dvss.n482 1.34003
R8069 dvss.n1628 dvss.n482 1.34003
R8070 dvss.n1274 dvss.n1273 1.34003
R8071 dvss.n1266 dvss.n1265 1.34003
R8072 dvss.n1265 dvss.n1264 1.34003
R8073 dvss.n1140 dvss.n601 1.34003
R8074 dvss.n1142 dvss.n592 1.34003
R8075 dvss.n1155 dvss.n592 1.34003
R8076 dvss.n790 dvss.n785 1.34003
R8077 dvss.n795 dvss.n793 1.34003
R8078 dvss.n798 dvss.n795 1.34003
R8079 dvss.n3644 dvss 1.23235
R8080 dvss.n67 dvss.n4 1.09487
R8081 dvss.n26 dvss.n25 1.05227
R8082 dvss.n67 dvss.n66 0.886661
R8083 dvss.n3525 dvss 0.856314
R8084 dvss.n3524 dvss.n3523 0.856314
R8085 dvss dvss.n3513 0.856314
R8086 dvss.n3280 dvss 0.856314
R8087 dvss.n3296 dvss.n245 0.856314
R8088 dvss.n3300 dvss 0.856314
R8089 dvss.n3162 dvss 0.856314
R8090 dvss.n3181 dvss.n310 0.856314
R8091 dvss.n3185 dvss 0.856314
R8092 dvss dvss.n3061 0.856314
R8093 dvss.n3069 dvss.n3062 0.856314
R8094 dvss.n3067 dvss 0.856314
R8095 dvss.n2937 dvss 0.856314
R8096 dvss.n2948 dvss.n432 0.856314
R8097 dvss.n2952 dvss 0.856314
R8098 dvss.n1559 dvss 0.856314
R8099 dvss.n1558 dvss.n1557 0.856314
R8100 dvss dvss.n1547 0.856314
R8101 dvss.n1345 dvss 0.856314
R8102 dvss.n1356 dvss.n541 0.856314
R8103 dvss.n1360 dvss 0.856314
R8104 dvss dvss.n1069 0.856314
R8105 dvss.n1072 dvss.n1070 0.856314
R8106 dvss dvss.n1076 0.856314
R8107 dvss dvss.n974 0.856314
R8108 dvss.n976 dvss.n975 0.856314
R8109 dvss dvss.n995 0.856314
R8110 dvss dvss.n3581 0.856314
R8111 dvss.n3583 dvss.n3582 0.856314
R8112 dvss dvss.n3597 0.856314
R8113 dvss.n2713 dvss 0.856314
R8114 dvss.n2706 dvss.n1762 0.856314
R8115 dvss.n2704 dvss 0.856314
R8116 dvss.n2763 dvss 0.856314
R8117 dvss.n2756 dvss.n1731 0.856314
R8118 dvss.n2754 dvss 0.856314
R8119 dvss.n2813 dvss 0.856314
R8120 dvss.n2806 dvss.n1700 0.856314
R8121 dvss.n2804 dvss 0.856314
R8122 dvss.n2863 dvss 0.856314
R8123 dvss.n2856 dvss.n1669 0.856314
R8124 dvss.n2854 dvss 0.856314
R8125 dvss dvss.n1613 0.856314
R8126 dvss.n1615 dvss.n1614 0.856314
R8127 dvss dvss.n1628 0.856314
R8128 dvss.n1273 dvss 0.856314
R8129 dvss.n1266 dvss.n1196 0.856314
R8130 dvss.n1264 dvss 0.856314
R8131 dvss dvss.n1140 0.856314
R8132 dvss.n1142 dvss.n1141 0.856314
R8133 dvss dvss.n1155 0.856314
R8134 dvss dvss.n790 0.856314
R8135 dvss.n793 dvss.n791 0.856314
R8136 dvss dvss.n798 0.856314
R8137 dvss.n60 dvss.n4 0.7755
R8138 dvss.n64 dvss.n63 0.7755
R8139 dvss.n66 dvss.n65 0.705857
R8140 dvss.n128 dvss.t117 0.627052
R8141 dvss.n126 dvss.t116 0.627052
R8142 dvss.n127 dvss.n126 0.5805
R8143 dvss.n129 dvss.n128 0.5805
R8144 dvss dvss.n3645 0.543548
R8145 dvss.n64 dvss.n8 0.529518
R8146 dvss.n51 dvss.n50 0.526527
R8147 dvss.n130 dvss.n127 0.279444
R8148 dvss.n130 dvss.n129 0.268206
R8149 dvss.n7 dvss.n4 0.2505
R8150 dvss.n878 dvss 0.215174
R8151 dvss.n879 dvss 0.215174
R8152 dvss.n884 dvss 0.215174
R8153 dvss dvss.n2663 0.215174
R8154 dvss dvss.n2662 0.215174
R8155 dvss.n2659 dvss 0.215174
R8156 dvss.n3742 dvss 0.187023
R8157 dvss.n65 dvss.n64 0.176839
R8158 dvss.n26 dvss.n21 0.120292
R8159 dvss.n33 dvss.n21 0.120292
R8160 dvss.n34 dvss.n33 0.120292
R8161 dvss.n35 dvss.n34 0.120292
R8162 dvss.n35 dvss.n18 0.120292
R8163 dvss.n42 dvss.n18 0.120292
R8164 dvss.n43 dvss.n42 0.120292
R8165 dvss.n54 dvss.n43 0.120292
R8166 dvss.n54 dvss.n53 0.120292
R8167 dvss.n53 dvss.n44 0.120292
R8168 dvss.n48 dvss.n44 0.120292
R8169 dvss.n48 dvss.n47 0.120292
R8170 dvss.n3751 dvss.n0 0.120292
R8171 dvss.n3746 dvss.n0 0.120292
R8172 dvss.n3746 dvss.n3745 0.120292
R8173 dvss.n3745 dvss.n3744 0.120292
R8174 dvss dvss.n2657 0.067223
R8175 dvss dvss.n2656 0.067223
R8176 dvss.n2653 dvss 0.067223
R8177 dvss dvss.n2652 0.067223
R8178 dvss dvss.n2651 0.067223
R8179 dvss.n2648 dvss 0.067223
R8180 dvss dvss.n2647 0.067223
R8181 dvss.n2640 dvss 0.067223
R8182 dvss dvss.n2639 0.067223
R8183 dvss.n2632 dvss 0.067223
R8184 dvss.n2628 dvss 0.067223
R8185 dvss.n2621 dvss 0.067223
R8186 dvss dvss.n2620 0.067223
R8187 dvss dvss.n2619 0.067223
R8188 dvss.n2616 dvss 0.067223
R8189 dvss dvss.n2615 0.067223
R8190 dvss dvss.n2614 0.067223
R8191 dvss.n2611 dvss 0.067223
R8192 dvss.n2603 dvss 0.067223
R8193 dvss.n2595 dvss 0.067223
R8194 dvss dvss.n2594 0.067223
R8195 dvss.n2587 dvss 0.067223
R8196 dvss dvss.n2586 0.067223
R8197 dvss dvss.n2585 0.067223
R8198 dvss dvss.n2581 0.067223
R8199 dvss.n2574 dvss 0.067223
R8200 dvss dvss.n2573 0.067223
R8201 dvss dvss.n2572 0.067223
R8202 dvss.n2569 dvss 0.067223
R8203 dvss dvss.n2568 0.067223
R8204 dvss dvss.n2567 0.067223
R8205 dvss.n2564 dvss 0.067223
R8206 dvss.n2556 dvss 0.067223
R8207 dvss.n2548 dvss 0.067223
R8208 dvss dvss.n2547 0.067223
R8209 dvss.n2540 dvss 0.067223
R8210 dvss dvss.n2539 0.067223
R8211 dvss dvss.n2538 0.067223
R8212 dvss dvss.n2534 0.067223
R8213 dvss.n2527 dvss 0.067223
R8214 dvss dvss.n2526 0.067223
R8215 dvss dvss.n2525 0.067223
R8216 dvss.n2522 dvss 0.067223
R8217 dvss dvss.n2521 0.067223
R8218 dvss dvss.n2520 0.067223
R8219 dvss.n2517 dvss 0.067223
R8220 dvss.n2509 dvss 0.067223
R8221 dvss.n2501 dvss 0.067223
R8222 dvss dvss.n2500 0.067223
R8223 dvss.n2493 dvss 0.067223
R8224 dvss dvss.n2492 0.067223
R8225 dvss dvss.n2491 0.067223
R8226 dvss dvss.n2487 0.067223
R8227 dvss.n2480 dvss 0.067223
R8228 dvss dvss.n2479 0.067223
R8229 dvss dvss.n2478 0.067223
R8230 dvss.n2475 dvss 0.067223
R8231 dvss dvss.n2474 0.067223
R8232 dvss dvss.n2473 0.067223
R8233 dvss.n2470 dvss 0.067223
R8234 dvss.n2462 dvss 0.067223
R8235 dvss.n2454 dvss 0.067223
R8236 dvss dvss.n2453 0.067223
R8237 dvss.n2446 dvss 0.067223
R8238 dvss dvss.n2445 0.067223
R8239 dvss dvss.n2444 0.067223
R8240 dvss dvss.n2440 0.067223
R8241 dvss.n2433 dvss 0.067223
R8242 dvss dvss.n2432 0.067223
R8243 dvss dvss.n2431 0.067223
R8244 dvss.n2428 dvss 0.067223
R8245 dvss dvss.n2427 0.067223
R8246 dvss dvss.n2426 0.067223
R8247 dvss.n2423 dvss 0.067223
R8248 dvss.n2415 dvss 0.067223
R8249 dvss.n2407 dvss 0.067223
R8250 dvss dvss.n2406 0.067223
R8251 dvss.n2399 dvss 0.067223
R8252 dvss dvss.n2398 0.067223
R8253 dvss dvss.n2397 0.067223
R8254 dvss dvss.n2393 0.067223
R8255 dvss.n2386 dvss 0.067223
R8256 dvss dvss.n2385 0.067223
R8257 dvss dvss.n2384 0.067223
R8258 dvss.n2381 dvss 0.067223
R8259 dvss dvss.n2380 0.067223
R8260 dvss dvss.n2379 0.067223
R8261 dvss.n2376 dvss 0.067223
R8262 dvss.n2368 dvss 0.067223
R8263 dvss.n2360 dvss 0.067223
R8264 dvss dvss.n2359 0.067223
R8265 dvss.n2352 dvss 0.067223
R8266 dvss dvss.n2351 0.067223
R8267 dvss dvss.n2350 0.067223
R8268 dvss dvss.n2346 0.067223
R8269 dvss.n2339 dvss 0.067223
R8270 dvss dvss.n2338 0.067223
R8271 dvss dvss.n2337 0.067223
R8272 dvss.n2334 dvss 0.067223
R8273 dvss dvss.n2333 0.067223
R8274 dvss dvss.n2332 0.067223
R8275 dvss.n2329 dvss 0.067223
R8276 dvss.n2321 dvss 0.067223
R8277 dvss.n2313 dvss 0.067223
R8278 dvss dvss.n2312 0.067223
R8279 dvss.n2305 dvss 0.067223
R8280 dvss dvss.n2304 0.067223
R8281 dvss dvss.n2303 0.067223
R8282 dvss dvss.n2299 0.067223
R8283 dvss.n3737 dvss 0.067223
R8284 dvss dvss.n3736 0.067223
R8285 dvss dvss.n3735 0.067223
R8286 dvss.n3732 dvss 0.067223
R8287 dvss dvss.n3731 0.067223
R8288 dvss dvss.n3730 0.067223
R8289 dvss.n3727 dvss 0.067223
R8290 dvss.n3719 dvss 0.067223
R8291 dvss.n3711 dvss 0.067223
R8292 dvss dvss.n3710 0.067223
R8293 dvss.n3703 dvss 0.067223
R8294 dvss dvss.n3702 0.067223
R8295 dvss dvss.n3701 0.067223
R8296 dvss dvss.n3697 0.067223
R8297 dvss.n3690 dvss 0.067223
R8298 dvss dvss.n3689 0.067223
R8299 dvss dvss.n3688 0.067223
R8300 dvss.n3685 dvss 0.067223
R8301 dvss dvss.n3684 0.067223
R8302 dvss dvss.n3683 0.067223
R8303 dvss.n3680 dvss 0.067223
R8304 dvss.n3672 dvss 0.067223
R8305 dvss.n3664 dvss 0.067223
R8306 dvss dvss.n3663 0.067223
R8307 dvss.n3656 dvss 0.067223
R8308 dvss dvss.n3655 0.067223
R8309 dvss dvss.n3654 0.067223
R8310 dvss dvss.n2602 0.0638446
R8311 dvss dvss.n2555 0.0638446
R8312 dvss dvss.n2508 0.0638446
R8313 dvss dvss.n2461 0.0638446
R8314 dvss dvss.n2414 0.0638446
R8315 dvss dvss.n2367 0.0638446
R8316 dvss dvss.n2320 0.0638446
R8317 dvss dvss.n3718 0.0638446
R8318 dvss dvss.n3671 0.0638446
R8319 dvss dvss.n2624 0.0613108
R8320 dvss dvss.n2577 0.0613108
R8321 dvss dvss.n2530 0.0613108
R8322 dvss dvss.n2483 0.0613108
R8323 dvss dvss.n2436 0.0613108
R8324 dvss dvss.n2389 0.0613108
R8325 dvss dvss.n2342 0.0613108
R8326 dvss dvss.n3693 0.0613108
R8327 dvss dvss.n3751 0.0603958
R8328 dvss.n3741 dvss 0.0520203
R8329 dvss.n129 dvss.t115 0.047052
R8330 dvss.n128 dvss.t119 0.047052
R8331 dvss.n126 dvss.t120 0.047052
R8332 dvss.n127 dvss.t118 0.047052
R8333 dvss.n2644 dvss 0.0469527
R8334 dvss.n2591 dvss 0.0469527
R8335 dvss.n2544 dvss 0.0469527
R8336 dvss.n2497 dvss 0.0469527
R8337 dvss.n2450 dvss 0.0469527
R8338 dvss.n2403 dvss 0.0469527
R8339 dvss.n2356 dvss 0.0469527
R8340 dvss.n2309 dvss 0.0469527
R8341 dvss.n3707 dvss 0.0469527
R8342 dvss.n3660 dvss 0.0469527
R8343 dvss dvss.n878 0.0466957
R8344 dvss dvss.n879 0.0466957
R8345 dvss.n2663 dvss 0.0466957
R8346 dvss.n2662 dvss 0.0466957
R8347 dvss dvss.n2610 0.0435743
R8348 dvss.n2599 dvss 0.0435743
R8349 dvss dvss.n2563 0.0435743
R8350 dvss.n2552 dvss 0.0435743
R8351 dvss dvss.n2516 0.0435743
R8352 dvss.n2505 dvss 0.0435743
R8353 dvss dvss.n2469 0.0435743
R8354 dvss.n2458 dvss 0.0435743
R8355 dvss dvss.n2422 0.0435743
R8356 dvss.n2411 dvss 0.0435743
R8357 dvss dvss.n2375 0.0435743
R8358 dvss.n2364 dvss 0.0435743
R8359 dvss dvss.n2328 0.0435743
R8360 dvss.n2317 dvss 0.0435743
R8361 dvss dvss.n3726 0.0435743
R8362 dvss.n3715 dvss 0.0435743
R8363 dvss dvss.n3679 0.0435743
R8364 dvss.n3668 dvss 0.0435743
R8365 dvss dvss.n2631 0.0410405
R8366 dvss.n2000 dvss 0.0410405
R8367 dvss.n2582 dvss 0.0410405
R8368 dvss.n2033 dvss 0.0410405
R8369 dvss.n2535 dvss 0.0410405
R8370 dvss.n2069 dvss 0.0410405
R8371 dvss.n2488 dvss 0.0410405
R8372 dvss.n2105 dvss 0.0410405
R8373 dvss.n2441 dvss 0.0410405
R8374 dvss.n2141 dvss 0.0410405
R8375 dvss.n2394 dvss 0.0410405
R8376 dvss.n2177 dvss 0.0410405
R8377 dvss.n2347 dvss 0.0410405
R8378 dvss.n2209 dvss 0.0410405
R8379 dvss.n2300 dvss 0.0410405
R8380 dvss.n2295 dvss 0.0410405
R8381 dvss.n3698 dvss 0.0410405
R8382 dvss.n95 dvss 0.0410405
R8383 dvss dvss.n2638 0.0385068
R8384 dvss.n885 dvss.n884 0.0358261
R8385 dvss.n2659 dvss.n2658 0.0358261
R8386 dvss dvss.n2635 0.0351284
R8387 dvss.n769 dvss 0.0323548
R8388 dvss.n770 dvss 0.0323548
R8389 dvss.n786 dvss 0.0323548
R8390 dvss.n777 dvss 0.0323548
R8391 dvss dvss.n782 0.0323548
R8392 dvss.n808 dvss 0.0323548
R8393 dvss.n809 dvss 0.0323548
R8394 dvss.n820 dvss 0.0323548
R8395 dvss dvss.n819 0.0323548
R8396 dvss.n1114 dvss 0.0323548
R8397 dvss.n1115 dvss 0.0323548
R8398 dvss.n1117 dvss 0.0323548
R8399 dvss dvss.n1116 0.0323548
R8400 dvss.n1126 dvss 0.0323548
R8401 dvss.n1129 dvss 0.0323548
R8402 dvss dvss.n1128 0.0323548
R8403 dvss.n1144 dvss 0.0323548
R8404 dvss dvss.n593 0.0323548
R8405 dvss.n1168 dvss 0.0323548
R8406 dvss.n1169 dvss 0.0323548
R8407 dvss.n1182 dvss 0.0323548
R8408 dvss.n1183 dvss 0.0323548
R8409 dvss.n1287 dvss 0.0323548
R8410 dvss dvss.n1286 0.0323548
R8411 dvss dvss.n1285 0.0323548
R8412 dvss.n1282 dvss 0.0323548
R8413 dvss dvss.n1280 0.0323548
R8414 dvss.n1277 dvss 0.0323548
R8415 dvss dvss.n1276 0.0323548
R8416 dvss.n1268 dvss 0.0323548
R8417 dvss.n1259 dvss 0.0323548
R8418 dvss.n1251 dvss 0.0323548
R8419 dvss dvss.n1250 0.0323548
R8420 dvss.n1241 dvss 0.0323548
R8421 dvss dvss.n1240 0.0323548
R8422 dvss.n1587 dvss 0.0323548
R8423 dvss.n1588 dvss 0.0323548
R8424 dvss.n1590 dvss 0.0323548
R8425 dvss dvss.n1589 0.0323548
R8426 dvss.n1599 dvss 0.0323548
R8427 dvss.n1602 dvss 0.0323548
R8428 dvss dvss.n1601 0.0323548
R8429 dvss.n1617 dvss 0.0323548
R8430 dvss dvss.n483 0.0323548
R8431 dvss.n1641 dvss 0.0323548
R8432 dvss.n1642 dvss 0.0323548
R8433 dvss.n1655 dvss 0.0323548
R8434 dvss.n1656 dvss 0.0323548
R8435 dvss.n2877 dvss 0.0323548
R8436 dvss dvss.n2876 0.0323548
R8437 dvss dvss.n2875 0.0323548
R8438 dvss.n2872 dvss 0.0323548
R8439 dvss dvss.n2870 0.0323548
R8440 dvss.n2867 dvss 0.0323548
R8441 dvss dvss.n2866 0.0323548
R8442 dvss.n2858 dvss 0.0323548
R8443 dvss.n2849 dvss 0.0323548
R8444 dvss.n2841 dvss 0.0323548
R8445 dvss dvss.n2840 0.0323548
R8446 dvss.n2831 dvss 0.0323548
R8447 dvss dvss.n2830 0.0323548
R8448 dvss dvss.n2829 0.0323548
R8449 dvss.n2826 dvss 0.0323548
R8450 dvss dvss.n2825 0.0323548
R8451 dvss dvss.n2824 0.0323548
R8452 dvss dvss.n2820 0.0323548
R8453 dvss dvss.n2819 0.0323548
R8454 dvss.n2816 dvss 0.0323548
R8455 dvss.n2808 dvss 0.0323548
R8456 dvss.n2799 dvss 0.0323548
R8457 dvss.n2791 dvss 0.0323548
R8458 dvss dvss.n2790 0.0323548
R8459 dvss.n2781 dvss 0.0323548
R8460 dvss dvss.n2780 0.0323548
R8461 dvss dvss.n2779 0.0323548
R8462 dvss.n2776 dvss 0.0323548
R8463 dvss dvss.n2775 0.0323548
R8464 dvss dvss.n2774 0.0323548
R8465 dvss dvss.n2770 0.0323548
R8466 dvss dvss.n2769 0.0323548
R8467 dvss.n2766 dvss 0.0323548
R8468 dvss.n2758 dvss 0.0323548
R8469 dvss.n2749 dvss 0.0323548
R8470 dvss.n2741 dvss 0.0323548
R8471 dvss dvss.n2740 0.0323548
R8472 dvss.n2731 dvss 0.0323548
R8473 dvss dvss.n2730 0.0323548
R8474 dvss dvss.n2729 0.0323548
R8475 dvss.n2726 dvss 0.0323548
R8476 dvss dvss.n2725 0.0323548
R8477 dvss dvss.n2724 0.0323548
R8478 dvss dvss.n2720 0.0323548
R8479 dvss dvss.n2719 0.0323548
R8480 dvss.n2716 dvss 0.0323548
R8481 dvss.n2708 dvss 0.0323548
R8482 dvss.n2699 dvss 0.0323548
R8483 dvss.n2691 dvss 0.0323548
R8484 dvss dvss.n2690 0.0323548
R8485 dvss dvss.n1775 0.0323548
R8486 dvss.n3552 dvss 0.0323548
R8487 dvss.n3553 dvss 0.0323548
R8488 dvss.n3567 dvss 0.0323548
R8489 dvss dvss.n3566 0.0323548
R8490 dvss dvss.n3565 0.0323548
R8491 dvss dvss.n3561 0.0323548
R8492 dvss dvss.n3560 0.0323548
R8493 dvss.n3577 dvss 0.0323548
R8494 dvss dvss.n3585 0.0323548
R8495 dvss.n3601 dvss 0.0323548
R8496 dvss.n3610 dvss 0.0323548
R8497 dvss.n3619 dvss 0.0323548
R8498 dvss.n3628 dvss 0.0323548
R8499 dvss.n3632 dvss 0.0323548
R8500 dvss dvss.n3631 0.0323548
R8501 dvss dvss.n3630 0.0323548
R8502 dvss dvss.n3629 0.0323548
R8503 dvss.n3643 dvss 0.0323548
R8504 dvss.n800 dvss 0.0319516
R8505 dvss dvss.n589 0.0319516
R8506 dvss dvss.n1258 0.0319516
R8507 dvss dvss.n479 0.0319516
R8508 dvss dvss.n2848 0.0319516
R8509 dvss dvss.n2798 0.0319516
R8510 dvss dvss.n2748 0.0319516
R8511 dvss dvss.n2698 0.0319516
R8512 dvss dvss.n3600 0.0319516
R8513 dvss dvss.n2606 0.0300608
R8514 dvss dvss.n2559 0.0300608
R8515 dvss dvss.n2512 0.0300608
R8516 dvss dvss.n2465 0.0300608
R8517 dvss dvss.n2418 0.0300608
R8518 dvss dvss.n2371 0.0300608
R8519 dvss dvss.n2324 0.0300608
R8520 dvss dvss.n3722 0.0300608
R8521 dvss dvss.n3675 0.0300608
R8522 dvss.n886 dvss 0.0282388
R8523 dvss.n888 dvss 0.0282388
R8524 dvss dvss.n887 0.0282388
R8525 dvss.n919 dvss 0.0282388
R8526 dvss dvss.n918 0.0282388
R8527 dvss.n929 dvss 0.0282388
R8528 dvss.n930 dvss 0.0282388
R8529 dvss dvss.n931 0.0282388
R8530 dvss.n955 dvss 0.0282388
R8531 dvss.n978 dvss 0.0282388
R8532 dvss.n984 dvss 0.0282388
R8533 dvss dvss.n1015 0.0282388
R8534 dvss dvss.n1029 0.0282388
R8535 dvss.n1040 dvss 0.0282388
R8536 dvss.n621 dvss 0.0282388
R8537 dvss.n622 dvss 0.0282388
R8538 dvss.n1049 dvss 0.0282388
R8539 dvss.n1058 dvss 0.0282388
R8540 dvss dvss.n640 0.0282388
R8541 dvss.n1080 dvss 0.0282388
R8542 dvss dvss.n703 0.0282388
R8543 dvss.n690 dvss 0.0282388
R8544 dvss.n1296 dvss 0.0282388
R8545 dvss dvss.n563 0.0282388
R8546 dvss.n1318 dvss 0.0282388
R8547 dvss.n1315 dvss 0.0282388
R8548 dvss.n1328 dvss 0.0282388
R8549 dvss.n1354 dvss 0.0282388
R8550 dvss dvss.n1365 0.0282388
R8551 dvss dvss.n1392 0.0282388
R8552 dvss dvss.n1406 0.0282388
R8553 dvss.n1416 dvss 0.0282388
R8554 dvss.n1574 dvss 0.0282388
R8555 dvss dvss.n1573 0.0282388
R8556 dvss dvss.n1572 0.0282388
R8557 dvss dvss.n1568 0.0282388
R8558 dvss.n1500 dvss 0.0282388
R8559 dvss dvss.n1551 0.0282388
R8560 dvss dvss.n1540 0.0282388
R8561 dvss.n1527 dvss 0.0282388
R8562 dvss.n2886 dvss 0.0282388
R8563 dvss.n2911 dvss 0.0282388
R8564 dvss.n2908 dvss 0.0282388
R8565 dvss dvss.n2907 0.0282388
R8566 dvss.n2920 dvss 0.0282388
R8567 dvss.n2946 dvss 0.0282388
R8568 dvss dvss.n2957 0.0282388
R8569 dvss dvss.n2984 0.0282388
R8570 dvss dvss.n2999 0.0282388
R8571 dvss.n3009 dvss 0.0282388
R8572 dvss dvss.n402 0.0282388
R8573 dvss.n3031 dvss 0.0282388
R8574 dvss.n3028 dvss 0.0282388
R8575 dvss.n3039 dvss 0.0282388
R8576 dvss.n3071 dvss 0.0282388
R8577 dvss.n3083 dvss 0.0282388
R8578 dvss.n3105 dvss 0.0282388
R8579 dvss dvss.n3116 0.0282388
R8580 dvss.n3126 dvss 0.0282388
R8581 dvss dvss.n3129 0.0282388
R8582 dvss.n3144 dvss 0.0282388
R8583 dvss dvss.n3143 0.0282388
R8584 dvss.n3153 dvss 0.0282388
R8585 dvss.n3179 dvss 0.0282388
R8586 dvss.n3199 dvss 0.0282388
R8587 dvss.n3221 dvss 0.0282388
R8588 dvss dvss.n3232 0.0282388
R8589 dvss.n3242 dvss 0.0282388
R8590 dvss dvss.n3245 0.0282388
R8591 dvss.n3260 dvss 0.0282388
R8592 dvss dvss.n3259 0.0282388
R8593 dvss.n3268 dvss 0.0282388
R8594 dvss.n3294 dvss 0.0282388
R8595 dvss dvss.n3302 0.0282388
R8596 dvss dvss.n3332 0.0282388
R8597 dvss dvss.n3346 0.0282388
R8598 dvss.n3356 dvss 0.0282388
R8599 dvss.n3540 dvss 0.0282388
R8600 dvss dvss.n3539 0.0282388
R8601 dvss dvss.n3538 0.0282388
R8602 dvss dvss.n3534 0.0282388
R8603 dvss.n3427 dvss 0.0282388
R8604 dvss dvss.n3517 0.0282388
R8605 dvss dvss.n3506 0.0282388
R8606 dvss dvss.n3418 0.0282388
R8607 dvss dvss.n3417 0.0282388
R8608 dvss.n3491 dvss 0.0282388
R8609 dvss dvss.n3490 0.0282388
R8610 dvss.n3646 dvss 0.0282388
R8611 dvss dvss.n742 0.0278876
R8612 dvss dvss.n1079 0.0278876
R8613 dvss.n1379 dvss 0.0278876
R8614 dvss dvss.n1550 0.0278876
R8615 dvss.n2971 dvss 0.0278876
R8616 dvss.n3087 dvss 0.0278876
R8617 dvss.n3203 dvss 0.0278876
R8618 dvss.n3319 dvss 0.0278876
R8619 dvss dvss.n3516 0.0278876
R8620 dvss.n963 dvss 0.0257809
R8621 dvss dvss.n632 0.0257809
R8622 dvss.n1334 dvss 0.0257809
R8623 dvss dvss.n1564 0.0257809
R8624 dvss.n2926 dvss 0.0257809
R8625 dvss.n3048 dvss 0.0257809
R8626 dvss.n3165 dvss 0.0257809
R8627 dvss.n3283 dvss 0.0257809
R8628 dvss dvss.n3530 0.0257809
R8629 dvss.n910 dvss 0.0250787
R8630 dvss.n2607 dvss 0.0233041
R8631 dvss.n2560 dvss 0.0233041
R8632 dvss.n2513 dvss 0.0233041
R8633 dvss.n2466 dvss 0.0233041
R8634 dvss.n2419 dvss 0.0233041
R8635 dvss.n2372 dvss 0.0233041
R8636 dvss.n2325 dvss 0.0233041
R8637 dvss.n3723 dvss 0.0233041
R8638 dvss.n3676 dvss 0.0233041
R8639 dvss dvss.n776 0.0230806
R8640 dvss dvss.n1138 0.0230806
R8641 dvss dvss.n1271 0.0230806
R8642 dvss dvss.n1611 0.0230806
R8643 dvss dvss.n2861 0.0230806
R8644 dvss dvss.n2811 0.0230806
R8645 dvss dvss.n2761 0.0230806
R8646 dvss dvss.n2711 0.0230806
R8647 dvss.n3586 dvss 0.0230806
R8648 dvss.n817 dvss 0.0226774
R8649 dvss.n583 dvss 0.0226774
R8650 dvss dvss.n1245 0.0226774
R8651 dvss.n473 dvss 0.0226774
R8652 dvss dvss.n2835 0.0226774
R8653 dvss dvss.n2785 0.0226774
R8654 dvss dvss.n2735 0.0226774
R8655 dvss dvss.n2685 0.0226774
R8656 dvss dvss.n3614 0.0226774
R8657 dvss.n47 dvss 0.0226354
R8658 dvss.n3744 dvss 0.0226354
R8659 dvss.n792 dvss 0.0222742
R8660 dvss.n802 dvss 0.0222742
R8661 dvss dvss.n1143 0.0222742
R8662 dvss dvss.n1158 0.0222742
R8663 dvss dvss.n1267 0.0222742
R8664 dvss.n1255 dvss 0.0222742
R8665 dvss dvss.n1616 0.0222742
R8666 dvss dvss.n1631 0.0222742
R8667 dvss dvss.n2857 0.0222742
R8668 dvss.n2845 dvss 0.0222742
R8669 dvss dvss.n2807 0.0222742
R8670 dvss.n2795 dvss 0.0222742
R8671 dvss dvss.n2757 0.0222742
R8672 dvss.n2745 dvss 0.0222742
R8673 dvss dvss.n2707 0.0222742
R8674 dvss.n2695 dvss 0.0222742
R8675 dvss dvss.n3584 0.0222742
R8676 dvss.n151 dvss 0.0222742
R8677 dvss dvss.n810 0.0202581
R8678 dvss.n1174 dvss 0.0202581
R8679 dvss.n1208 dvss 0.0202581
R8680 dvss.n1647 dvss 0.0202581
R8681 dvss.n1681 dvss 0.0202581
R8682 dvss.n1712 dvss 0.0202581
R8683 dvss.n1743 dvss 0.0202581
R8684 dvss.n1774 dvss 0.0202581
R8685 dvss.n3613 dvss 0.0202581
R8686 dvss dvss.n972 0.0201629
R8687 dvss dvss.n1067 0.0201629
R8688 dvss.n1347 dvss 0.0201629
R8689 dvss.n1499 dvss 0.0201629
R8690 dvss.n2939 dvss 0.0201629
R8691 dvss dvss.n3059 0.0201629
R8692 dvss.n3176 dvss 0.0201629
R8693 dvss.n3293 dvss 0.0201629
R8694 dvss.n3426 dvss 0.0201629
R8695 dvss.n1125 dvss 0.0198548
R8696 dvss dvss.n1281 0.0198548
R8697 dvss.n1598 dvss 0.0198548
R8698 dvss dvss.n2871 0.0198548
R8699 dvss.n2821 dvss 0.0198548
R8700 dvss.n2771 dvss 0.0198548
R8701 dvss.n2721 dvss 0.0198548
R8702 dvss.n3562 dvss 0.0198548
R8703 dvss dvss.n868 0.0198118
R8704 dvss.n1037 dvss 0.0198118
R8705 dvss.n1299 dvss 0.0198118
R8706 dvss dvss.n511 0.0198118
R8707 dvss.n2889 dvss 0.0198118
R8708 dvss dvss.n401 0.0198118
R8709 dvss dvss.n339 0.0198118
R8710 dvss dvss.n275 0.0198118
R8711 dvss dvss.n212 0.0198118
R8712 dvss.n3495 dvss 0.0198118
R8713 dvss dvss.n977 0.0194607
R8714 dvss.n1071 dvss 0.0194607
R8715 dvss.n1355 dvss 0.0194607
R8716 dvss.n1556 dvss 0.0194607
R8717 dvss.n2947 dvss 0.0194607
R8718 dvss dvss.n3070 0.0194607
R8719 dvss.n3180 dvss 0.0194607
R8720 dvss.n3295 dvss 0.0194607
R8721 dvss.n3522 dvss 0.0194607
R8722 dvss dvss.n999 0.0184073
R8723 dvss.n652 dvss 0.0184073
R8724 dvss dvss.n532 0.0184073
R8725 dvss.n1449 dvss 0.0184073
R8726 dvss dvss.n423 0.0184073
R8727 dvss dvss.n363 0.0184073
R8728 dvss dvss.n299 0.0184073
R8729 dvss dvss.n233 0.0184073
R8730 dvss.n3389 dvss 0.0184073
R8731 dvss.n2636 dvss 0.0182365
R8732 dvss.n949 dvss 0.0173539
R8733 dvss dvss.n763 0.0173539
R8734 dvss.n1052 dvss 0.0173539
R8735 dvss dvss.n631 0.0173539
R8736 dvss dvss.n1314 0.0173539
R8737 dvss dvss.n552 0.0173539
R8738 dvss.n1569 dvss 0.0173539
R8739 dvss.n1429 dvss 0.0173539
R8740 dvss dvss.n2906 0.0173539
R8741 dvss dvss.n443 0.0173539
R8742 dvss dvss.n3027 0.0173539
R8743 dvss.n3045 dvss 0.0173539
R8744 dvss dvss.n3142 0.0173539
R8745 dvss dvss.n319 0.0173539
R8746 dvss dvss.n3258 0.0173539
R8747 dvss.n3274 dvss 0.0173539
R8748 dvss.n3535 dvss 0.0173539
R8749 dvss.n3369 dvss 0.0173539
R8750 dvss.n912 dvss 0.0166517
R8751 dvss.n934 dvss 0.0163006
R8752 dvss.n1034 dvss 0.0163006
R8753 dvss dvss.n722 0.0163006
R8754 dvss.n696 dvss 0.0163006
R8755 dvss dvss.n698 0.0163006
R8756 dvss.n1411 dvss 0.0163006
R8757 dvss dvss.n516 0.0163006
R8758 dvss.n1533 dvss 0.0163006
R8759 dvss dvss.n1535 0.0163006
R8760 dvss.n3004 dvss 0.0163006
R8761 dvss dvss.n407 0.0163006
R8762 dvss.n3121 dvss 0.0163006
R8763 dvss dvss.n344 0.0163006
R8764 dvss.n3237 dvss 0.0163006
R8765 dvss dvss.n280 0.0163006
R8766 dvss.n3351 dvss 0.0163006
R8767 dvss dvss.n217 0.0163006
R8768 dvss.n3499 dvss 0.0163006
R8769 dvss dvss.n3501 0.0163006
R8770 dvss dvss.n932 0.0148961
R8771 dvss.n2657 dvss 0.0148581
R8772 dvss.n2656 dvss 0.0148581
R8773 dvss.n2653 dvss 0.0148581
R8774 dvss.n2652 dvss 0.0148581
R8775 dvss.n2651 dvss 0.0148581
R8776 dvss.n2648 dvss 0.0148581
R8777 dvss.n2647 dvss 0.0148581
R8778 dvss.n2646 dvss 0.0148581
R8779 dvss.n2640 dvss 0.0148581
R8780 dvss.n2639 dvss 0.0148581
R8781 dvss.n2638 dvss 0.0148581
R8782 dvss.n1989 dvss 0.0148581
R8783 dvss.n1989 dvss 0.0148581
R8784 dvss.n2636 dvss 0.0148581
R8785 dvss.n2635 dvss 0.0148581
R8786 dvss.n2632 dvss 0.0148581
R8787 dvss.n2631 dvss 0.0148581
R8788 dvss.n2628 dvss 0.0148581
R8789 dvss.n2627 dvss 0.0148581
R8790 dvss.n2624 dvss 0.0148581
R8791 dvss.n2621 dvss 0.0148581
R8792 dvss.n2620 dvss 0.0148581
R8793 dvss.n2619 dvss 0.0148581
R8794 dvss.n2616 dvss 0.0148581
R8795 dvss.n2615 dvss 0.0148581
R8796 dvss.n2614 dvss 0.0148581
R8797 dvss.n2611 dvss 0.0148581
R8798 dvss.n2610 dvss 0.0148581
R8799 dvss dvss.n2013 0.0148581
R8800 dvss.n2607 dvss 0.0148581
R8801 dvss.n2606 dvss 0.0148581
R8802 dvss.n2603 dvss 0.0148581
R8803 dvss.n2599 dvss 0.0148581
R8804 dvss.n2598 dvss 0.0148581
R8805 dvss.n2595 dvss 0.0148581
R8806 dvss.n2594 dvss 0.0148581
R8807 dvss.n2593 dvss 0.0148581
R8808 dvss.n2587 dvss 0.0148581
R8809 dvss.n2586 dvss 0.0148581
R8810 dvss.n2585 dvss 0.0148581
R8811 dvss.n2582 dvss 0.0148581
R8812 dvss.n2581 dvss 0.0148581
R8813 dvss.n2580 dvss 0.0148581
R8814 dvss.n2577 dvss 0.0148581
R8815 dvss.n2574 dvss 0.0148581
R8816 dvss.n2573 dvss 0.0148581
R8817 dvss.n2572 dvss 0.0148581
R8818 dvss.n2569 dvss 0.0148581
R8819 dvss.n2568 dvss 0.0148581
R8820 dvss.n2567 dvss 0.0148581
R8821 dvss.n2564 dvss 0.0148581
R8822 dvss.n2563 dvss 0.0148581
R8823 dvss dvss.n2049 0.0148581
R8824 dvss.n2560 dvss 0.0148581
R8825 dvss.n2559 dvss 0.0148581
R8826 dvss.n2556 dvss 0.0148581
R8827 dvss.n2552 dvss 0.0148581
R8828 dvss.n2551 dvss 0.0148581
R8829 dvss.n2548 dvss 0.0148581
R8830 dvss.n2547 dvss 0.0148581
R8831 dvss.n2546 dvss 0.0148581
R8832 dvss.n2540 dvss 0.0148581
R8833 dvss.n2539 dvss 0.0148581
R8834 dvss.n2538 dvss 0.0148581
R8835 dvss.n2535 dvss 0.0148581
R8836 dvss.n2534 dvss 0.0148581
R8837 dvss.n2533 dvss 0.0148581
R8838 dvss.n2530 dvss 0.0148581
R8839 dvss.n2527 dvss 0.0148581
R8840 dvss.n2526 dvss 0.0148581
R8841 dvss.n2525 dvss 0.0148581
R8842 dvss.n2522 dvss 0.0148581
R8843 dvss.n2521 dvss 0.0148581
R8844 dvss.n2520 dvss 0.0148581
R8845 dvss.n2517 dvss 0.0148581
R8846 dvss.n2516 dvss 0.0148581
R8847 dvss dvss.n2085 0.0148581
R8848 dvss.n2513 dvss 0.0148581
R8849 dvss.n2512 dvss 0.0148581
R8850 dvss.n2509 dvss 0.0148581
R8851 dvss.n2505 dvss 0.0148581
R8852 dvss.n2504 dvss 0.0148581
R8853 dvss.n2501 dvss 0.0148581
R8854 dvss.n2500 dvss 0.0148581
R8855 dvss.n2499 dvss 0.0148581
R8856 dvss.n2493 dvss 0.0148581
R8857 dvss.n2492 dvss 0.0148581
R8858 dvss.n2491 dvss 0.0148581
R8859 dvss.n2488 dvss 0.0148581
R8860 dvss.n2487 dvss 0.0148581
R8861 dvss.n2486 dvss 0.0148581
R8862 dvss.n2483 dvss 0.0148581
R8863 dvss.n2480 dvss 0.0148581
R8864 dvss.n2479 dvss 0.0148581
R8865 dvss.n2478 dvss 0.0148581
R8866 dvss.n2475 dvss 0.0148581
R8867 dvss.n2474 dvss 0.0148581
R8868 dvss.n2473 dvss 0.0148581
R8869 dvss.n2470 dvss 0.0148581
R8870 dvss.n2469 dvss 0.0148581
R8871 dvss dvss.n2121 0.0148581
R8872 dvss.n2466 dvss 0.0148581
R8873 dvss.n2465 dvss 0.0148581
R8874 dvss.n2462 dvss 0.0148581
R8875 dvss.n2458 dvss 0.0148581
R8876 dvss.n2457 dvss 0.0148581
R8877 dvss.n2454 dvss 0.0148581
R8878 dvss.n2453 dvss 0.0148581
R8879 dvss.n2452 dvss 0.0148581
R8880 dvss.n2446 dvss 0.0148581
R8881 dvss.n2445 dvss 0.0148581
R8882 dvss.n2444 dvss 0.0148581
R8883 dvss.n2441 dvss 0.0148581
R8884 dvss.n2440 dvss 0.0148581
R8885 dvss.n2439 dvss 0.0148581
R8886 dvss.n2436 dvss 0.0148581
R8887 dvss.n2433 dvss 0.0148581
R8888 dvss.n2432 dvss 0.0148581
R8889 dvss.n2431 dvss 0.0148581
R8890 dvss.n2428 dvss 0.0148581
R8891 dvss.n2427 dvss 0.0148581
R8892 dvss.n2426 dvss 0.0148581
R8893 dvss.n2423 dvss 0.0148581
R8894 dvss.n2422 dvss 0.0148581
R8895 dvss dvss.n2157 0.0148581
R8896 dvss.n2419 dvss 0.0148581
R8897 dvss.n2418 dvss 0.0148581
R8898 dvss.n2415 dvss 0.0148581
R8899 dvss.n2411 dvss 0.0148581
R8900 dvss.n2410 dvss 0.0148581
R8901 dvss.n2407 dvss 0.0148581
R8902 dvss.n2406 dvss 0.0148581
R8903 dvss.n2405 dvss 0.0148581
R8904 dvss.n2399 dvss 0.0148581
R8905 dvss.n2398 dvss 0.0148581
R8906 dvss.n2397 dvss 0.0148581
R8907 dvss.n2394 dvss 0.0148581
R8908 dvss.n2393 dvss 0.0148581
R8909 dvss.n2392 dvss 0.0148581
R8910 dvss.n2389 dvss 0.0148581
R8911 dvss.n2386 dvss 0.0148581
R8912 dvss.n2385 dvss 0.0148581
R8913 dvss.n2384 dvss 0.0148581
R8914 dvss.n2381 dvss 0.0148581
R8915 dvss.n2380 dvss 0.0148581
R8916 dvss.n2379 dvss 0.0148581
R8917 dvss.n2376 dvss 0.0148581
R8918 dvss.n2375 dvss 0.0148581
R8919 dvss dvss.n2194 0.0148581
R8920 dvss.n2372 dvss 0.0148581
R8921 dvss.n2371 dvss 0.0148581
R8922 dvss.n2368 dvss 0.0148581
R8923 dvss.n2364 dvss 0.0148581
R8924 dvss.n2363 dvss 0.0148581
R8925 dvss.n2360 dvss 0.0148581
R8926 dvss.n2359 dvss 0.0148581
R8927 dvss.n2358 dvss 0.0148581
R8928 dvss.n2352 dvss 0.0148581
R8929 dvss.n2351 dvss 0.0148581
R8930 dvss.n2350 dvss 0.0148581
R8931 dvss.n2347 dvss 0.0148581
R8932 dvss.n2346 dvss 0.0148581
R8933 dvss.n2345 dvss 0.0148581
R8934 dvss.n2342 dvss 0.0148581
R8935 dvss.n2339 dvss 0.0148581
R8936 dvss.n2338 dvss 0.0148581
R8937 dvss.n2337 dvss 0.0148581
R8938 dvss.n2334 dvss 0.0148581
R8939 dvss.n2333 dvss 0.0148581
R8940 dvss.n2332 dvss 0.0148581
R8941 dvss.n2329 dvss 0.0148581
R8942 dvss.n2328 dvss 0.0148581
R8943 dvss dvss.n2248 0.0148581
R8944 dvss.n2325 dvss 0.0148581
R8945 dvss.n2324 dvss 0.0148581
R8946 dvss.n2321 dvss 0.0148581
R8947 dvss.n2317 dvss 0.0148581
R8948 dvss.n2316 dvss 0.0148581
R8949 dvss.n2313 dvss 0.0148581
R8950 dvss.n2312 dvss 0.0148581
R8951 dvss.n2311 dvss 0.0148581
R8952 dvss.n2305 dvss 0.0148581
R8953 dvss.n2304 dvss 0.0148581
R8954 dvss.n2303 dvss 0.0148581
R8955 dvss.n2300 dvss 0.0148581
R8956 dvss.n2299 dvss 0.0148581
R8957 dvss.n2298 dvss 0.0148581
R8958 dvss.n3740 dvss 0.0148581
R8959 dvss.n3737 dvss 0.0148581
R8960 dvss.n3736 dvss 0.0148581
R8961 dvss.n3735 dvss 0.0148581
R8962 dvss.n3732 dvss 0.0148581
R8963 dvss.n3731 dvss 0.0148581
R8964 dvss.n3730 dvss 0.0148581
R8965 dvss.n3727 dvss 0.0148581
R8966 dvss.n3726 dvss 0.0148581
R8967 dvss dvss.n79 0.0148581
R8968 dvss.n3723 dvss 0.0148581
R8969 dvss.n3722 dvss 0.0148581
R8970 dvss.n3719 dvss 0.0148581
R8971 dvss.n3715 dvss 0.0148581
R8972 dvss.n3714 dvss 0.0148581
R8973 dvss.n3711 dvss 0.0148581
R8974 dvss.n3710 dvss 0.0148581
R8975 dvss.n3709 dvss 0.0148581
R8976 dvss.n3703 dvss 0.0148581
R8977 dvss.n3702 dvss 0.0148581
R8978 dvss.n3701 dvss 0.0148581
R8979 dvss.n3698 dvss 0.0148581
R8980 dvss.n3697 dvss 0.0148581
R8981 dvss.n3696 dvss 0.0148581
R8982 dvss.n3693 dvss 0.0148581
R8983 dvss.n3690 dvss 0.0148581
R8984 dvss.n3689 dvss 0.0148581
R8985 dvss.n3688 dvss 0.0148581
R8986 dvss.n3685 dvss 0.0148581
R8987 dvss.n3684 dvss 0.0148581
R8988 dvss.n3683 dvss 0.0148581
R8989 dvss.n3680 dvss 0.0148581
R8990 dvss.n3679 dvss 0.0148581
R8991 dvss dvss.n107 0.0148581
R8992 dvss.n3676 dvss 0.0148581
R8993 dvss.n3675 dvss 0.0148581
R8994 dvss.n3672 dvss 0.0148581
R8995 dvss.n3668 dvss 0.0148581
R8996 dvss.n3667 dvss 0.0148581
R8997 dvss.n3664 dvss 0.0148581
R8998 dvss.n3663 dvss 0.0148581
R8999 dvss.n3662 dvss 0.0148581
R9000 dvss.n3656 dvss 0.0148581
R9001 dvss.n3655 dvss 0.0148581
R9002 dvss.n3654 dvss 0.0148581
R9003 dvss.n2643 dvss 0.0140135
R9004 dvss.n788 dvss 0.0134032
R9005 dvss dvss.n796 0.0134032
R9006 dvss.n1137 dvss 0.0134032
R9007 dvss dvss.n1153 0.0134032
R9008 dvss.n1191 dvss 0.0134032
R9009 dvss dvss.n1262 0.0134032
R9010 dvss.n1610 dvss 0.0134032
R9011 dvss dvss.n1626 0.0134032
R9012 dvss.n1664 dvss 0.0134032
R9013 dvss dvss.n2852 0.0134032
R9014 dvss.n1696 dvss 0.0134032
R9015 dvss dvss.n2802 0.0134032
R9016 dvss.n1727 dvss 0.0134032
R9017 dvss dvss.n2752 0.0134032
R9018 dvss.n1758 dvss 0.0134032
R9019 dvss dvss.n2702 0.0134032
R9020 dvss.n3579 dvss 0.0134032
R9021 dvss dvss.n3595 0.0134032
R9022 dvss.n768 dvss.n767 0.013
R9023 dvss.n1016 dvss 0.0127893
R9024 dvss.n704 dvss 0.0127893
R9025 dvss.n1393 dvss 0.0127893
R9026 dvss.n1541 dvss 0.0127893
R9027 dvss.n2985 dvss 0.0127893
R9028 dvss.n3098 dvss 0.0127893
R9029 dvss.n3214 dvss 0.0127893
R9030 dvss.n3333 dvss 0.0127893
R9031 dvss.n3507 dvss 0.0127893
R9032 dvss.n787 dvss 0.0125968
R9033 dvss.n797 dvss 0.0125968
R9034 dvss dvss.n1127 0.0125968
R9035 dvss.n1154 dvss 0.0125968
R9036 dvss dvss.n1275 0.0125968
R9037 dvss.n1263 dvss 0.0125968
R9038 dvss dvss.n1600 0.0125968
R9039 dvss.n1627 dvss 0.0125968
R9040 dvss dvss.n2865 0.0125968
R9041 dvss.n2853 dvss 0.0125968
R9042 dvss dvss.n2815 0.0125968
R9043 dvss.n2803 dvss 0.0125968
R9044 dvss dvss.n2765 0.0125968
R9045 dvss.n2753 dvss 0.0125968
R9046 dvss dvss.n2715 0.0125968
R9047 dvss.n2703 dvss 0.0125968
R9048 dvss.n3578 dvss 0.0125968
R9049 dvss.n3596 dvss 0.0125968
R9050 dvss dvss.n2627 0.0123243
R9051 dvss dvss.n2580 0.0123243
R9052 dvss dvss.n2533 0.0123243
R9053 dvss dvss.n2486 0.0123243
R9054 dvss dvss.n2439 0.0123243
R9055 dvss dvss.n2392 0.0123243
R9056 dvss dvss.n2345 0.0123243
R9057 dvss dvss.n2298 0.0123243
R9058 dvss dvss.n3696 0.0123243
R9059 dvss.n965 dvss 0.011736
R9060 dvss dvss.n993 0.011736
R9061 dvss dvss.n633 0.011736
R9062 dvss dvss.n642 0.011736
R9063 dvss dvss.n1341 0.011736
R9064 dvss.n1366 dvss 0.011736
R9065 dvss.n1561 dvss 0.011736
R9066 dvss.n1552 dvss 0.011736
R9067 dvss dvss.n2933 0.011736
R9068 dvss.n2958 dvss 0.011736
R9069 dvss dvss.n384 0.011736
R9070 dvss dvss.n3065 0.011736
R9071 dvss.n3160 dvss 0.011736
R9072 dvss dvss.n309 0.011736
R9073 dvss.n3278 dvss 0.011736
R9074 dvss.n3303 dvss 0.011736
R9075 dvss.n3527 dvss 0.011736
R9076 dvss.n3518 dvss 0.011736
R9077 dvss dvss.n2019 0.0114797
R9078 dvss.n2590 dvss 0.0114797
R9079 dvss dvss.n2055 0.0114797
R9080 dvss.n2543 dvss 0.0114797
R9081 dvss dvss.n2091 0.0114797
R9082 dvss.n2496 dvss 0.0114797
R9083 dvss dvss.n2127 0.0114797
R9084 dvss.n2449 dvss 0.0114797
R9085 dvss dvss.n2163 0.0114797
R9086 dvss.n2402 dvss 0.0114797
R9087 dvss dvss.n2197 0.0114797
R9088 dvss.n2355 dvss 0.0114797
R9089 dvss dvss.n2252 0.0114797
R9090 dvss.n2308 dvss 0.0114797
R9091 dvss dvss.n83 0.0114797
R9092 dvss.n3706 dvss 0.0114797
R9093 dvss dvss.n111 0.0114797
R9094 dvss.n3659 dvss 0.0114797
R9095 dvss.n885 dvss 0.0113696
R9096 dvss.n2658 dvss 0.0113696
R9097 dvss.n964 dvss 0.0110337
R9098 dvss.n994 dvss 0.0110337
R9099 dvss.n709 dvss 0.0110337
R9100 dvss.n1075 dvss 0.0110337
R9101 dvss.n1342 dvss 0.0110337
R9102 dvss dvss.n1361 0.0110337
R9103 dvss.n1436 dvss 0.0110337
R9104 dvss.n1546 dvss 0.0110337
R9105 dvss.n2934 dvss 0.0110337
R9106 dvss dvss.n2953 0.0110337
R9107 dvss dvss.n385 0.0110337
R9108 dvss.n3066 dvss 0.0110337
R9109 dvss dvss.n3164 0.0110337
R9110 dvss dvss.n3186 0.0110337
R9111 dvss dvss.n3282 0.0110337
R9112 dvss.n3301 dvss 0.0110337
R9113 dvss.n3376 dvss 0.0110337
R9114 dvss.n3512 dvss 0.0110337
R9115 dvss dvss.n737 0.00998034
R9116 dvss.n659 dvss 0.00998034
R9117 dvss dvss.n1382 0.00998034
R9118 dvss.n1457 dvss 0.00998034
R9119 dvss dvss.n2974 0.00998034
R9120 dvss dvss.n3090 0.00998034
R9121 dvss dvss.n3206 0.00998034
R9122 dvss dvss.n3322 0.00998034
R9123 dvss.n3401 dvss 0.00998034
R9124 dvss.n2013 dvss 0.00979054
R9125 dvss dvss.n2598 0.00979054
R9126 dvss.n2049 dvss 0.00979054
R9127 dvss dvss.n2551 0.00979054
R9128 dvss.n2085 dvss 0.00979054
R9129 dvss dvss.n2504 0.00979054
R9130 dvss.n2121 dvss 0.00979054
R9131 dvss dvss.n2457 0.00979054
R9132 dvss.n2157 dvss 0.00979054
R9133 dvss dvss.n2410 0.00979054
R9134 dvss.n2194 dvss 0.00979054
R9135 dvss dvss.n2363 0.00979054
R9136 dvss.n2248 dvss 0.00979054
R9137 dvss dvss.n2316 0.00979054
R9138 dvss.n3741 dvss.n3740 0.00979054
R9139 dvss.n79 dvss 0.00979054
R9140 dvss dvss.n3714 0.00979054
R9141 dvss.n107 dvss 0.00979054
R9142 dvss dvss.n3667 0.00979054
R9143 dvss.n2625 dvss 0.00894595
R9144 dvss.n2578 dvss 0.00894595
R9145 dvss.n2531 dvss 0.00894595
R9146 dvss.n2484 dvss 0.00894595
R9147 dvss.n2437 dvss 0.00894595
R9148 dvss.n2390 dvss 0.00894595
R9149 dvss.n2343 dvss 0.00894595
R9150 dvss.n2296 dvss 0.00894595
R9151 dvss.n3694 dvss 0.00894595
R9152 dvss dvss.n936 0.0078736
R9153 dvss dvss.n768 0.00735484
R9154 dvss dvss.n769 0.00735484
R9155 dvss dvss.n770 0.00735484
R9156 dvss dvss.n786 0.00735484
R9157 dvss dvss.n787 0.00735484
R9158 dvss dvss.n788 0.00735484
R9159 dvss.n789 dvss 0.00735484
R9160 dvss dvss.n776 0.00735484
R9161 dvss dvss.n777 0.00735484
R9162 dvss.n792 dvss 0.00735484
R9163 dvss dvss.n778 0.00735484
R9164 dvss.n797 dvss 0.00735484
R9165 dvss.n796 dvss 0.00735484
R9166 dvss dvss.n782 0.00735484
R9167 dvss dvss.n802 0.00735484
R9168 dvss dvss.n803 0.00735484
R9169 dvss dvss.n808 0.00735484
R9170 dvss dvss.n809 0.00735484
R9171 dvss.n811 dvss 0.00735484
R9172 dvss dvss.n817 0.00735484
R9173 dvss dvss.n818 0.00735484
R9174 dvss.n820 dvss 0.00735484
R9175 dvss.n819 dvss 0.00735484
R9176 dvss dvss.n1114 0.00735484
R9177 dvss dvss.n1115 0.00735484
R9178 dvss.n1117 dvss 0.00735484
R9179 dvss.n1116 dvss 0.00735484
R9180 dvss dvss.n1125 0.00735484
R9181 dvss dvss.n1126 0.00735484
R9182 dvss.n1129 dvss 0.00735484
R9183 dvss.n1128 dvss 0.00735484
R9184 dvss.n1127 dvss 0.00735484
R9185 dvss dvss.n1137 0.00735484
R9186 dvss.n1139 dvss 0.00735484
R9187 dvss.n1138 dvss 0.00735484
R9188 dvss.n1144 dvss 0.00735484
R9189 dvss.n1143 dvss 0.00735484
R9190 dvss.n599 dvss 0.00735484
R9191 dvss.n1154 dvss 0.00735484
R9192 dvss.n1153 dvss 0.00735484
R9193 dvss.n593 dvss 0.00735484
R9194 dvss.n1158 dvss 0.00735484
R9195 dvss.n590 dvss 0.00735484
R9196 dvss dvss.n1168 0.00735484
R9197 dvss dvss.n1169 0.00735484
R9198 dvss.n1170 dvss 0.00735484
R9199 dvss.n583 dvss 0.00735484
R9200 dvss.n582 dvss 0.00735484
R9201 dvss dvss.n1182 0.00735484
R9202 dvss dvss.n1183 0.00735484
R9203 dvss.n1287 dvss 0.00735484
R9204 dvss.n1286 dvss 0.00735484
R9205 dvss.n1285 dvss 0.00735484
R9206 dvss.n1282 dvss 0.00735484
R9207 dvss.n1281 dvss 0.00735484
R9208 dvss.n1280 dvss 0.00735484
R9209 dvss.n1277 dvss 0.00735484
R9210 dvss.n1276 dvss 0.00735484
R9211 dvss.n1275 dvss 0.00735484
R9212 dvss.n1191 dvss 0.00735484
R9213 dvss.n1272 dvss 0.00735484
R9214 dvss.n1271 dvss 0.00735484
R9215 dvss.n1268 dvss 0.00735484
R9216 dvss.n1267 dvss 0.00735484
R9217 dvss dvss.n1198 0.00735484
R9218 dvss.n1263 dvss 0.00735484
R9219 dvss.n1262 dvss 0.00735484
R9220 dvss.n1259 dvss 0.00735484
R9221 dvss.n1255 dvss 0.00735484
R9222 dvss.n1254 dvss 0.00735484
R9223 dvss.n1251 dvss 0.00735484
R9224 dvss.n1250 dvss 0.00735484
R9225 dvss.n1249 dvss 0.00735484
R9226 dvss.n1245 dvss 0.00735484
R9227 dvss.n1244 dvss 0.00735484
R9228 dvss.n1241 dvss 0.00735484
R9229 dvss.n1240 dvss 0.00735484
R9230 dvss dvss.n1587 0.00735484
R9231 dvss dvss.n1588 0.00735484
R9232 dvss.n1590 dvss 0.00735484
R9233 dvss.n1589 dvss 0.00735484
R9234 dvss dvss.n1598 0.00735484
R9235 dvss dvss.n1599 0.00735484
R9236 dvss.n1602 dvss 0.00735484
R9237 dvss.n1601 dvss 0.00735484
R9238 dvss.n1600 dvss 0.00735484
R9239 dvss dvss.n1610 0.00735484
R9240 dvss.n1612 dvss 0.00735484
R9241 dvss.n1611 dvss 0.00735484
R9242 dvss.n1617 dvss 0.00735484
R9243 dvss.n1616 dvss 0.00735484
R9244 dvss.n489 dvss 0.00735484
R9245 dvss.n1627 dvss 0.00735484
R9246 dvss.n1626 dvss 0.00735484
R9247 dvss.n483 dvss 0.00735484
R9248 dvss.n1631 dvss 0.00735484
R9249 dvss.n480 dvss 0.00735484
R9250 dvss dvss.n1641 0.00735484
R9251 dvss dvss.n1642 0.00735484
R9252 dvss.n1643 dvss 0.00735484
R9253 dvss.n473 dvss 0.00735484
R9254 dvss.n472 dvss 0.00735484
R9255 dvss dvss.n1655 0.00735484
R9256 dvss dvss.n1656 0.00735484
R9257 dvss.n2877 dvss 0.00735484
R9258 dvss.n2876 dvss 0.00735484
R9259 dvss.n2875 dvss 0.00735484
R9260 dvss.n2872 dvss 0.00735484
R9261 dvss.n2871 dvss 0.00735484
R9262 dvss.n2870 dvss 0.00735484
R9263 dvss.n2867 dvss 0.00735484
R9264 dvss.n2866 dvss 0.00735484
R9265 dvss.n2865 dvss 0.00735484
R9266 dvss.n1664 dvss 0.00735484
R9267 dvss.n2862 dvss 0.00735484
R9268 dvss.n2861 dvss 0.00735484
R9269 dvss.n2858 dvss 0.00735484
R9270 dvss.n2857 dvss 0.00735484
R9271 dvss dvss.n1671 0.00735484
R9272 dvss.n2853 dvss 0.00735484
R9273 dvss.n2852 dvss 0.00735484
R9274 dvss.n2849 dvss 0.00735484
R9275 dvss.n2845 dvss 0.00735484
R9276 dvss.n2844 dvss 0.00735484
R9277 dvss.n2841 dvss 0.00735484
R9278 dvss.n2840 dvss 0.00735484
R9279 dvss.n2839 dvss 0.00735484
R9280 dvss.n2835 dvss 0.00735484
R9281 dvss.n2834 dvss 0.00735484
R9282 dvss.n2831 dvss 0.00735484
R9283 dvss.n2830 dvss 0.00735484
R9284 dvss.n2829 dvss 0.00735484
R9285 dvss.n2826 dvss 0.00735484
R9286 dvss.n2825 dvss 0.00735484
R9287 dvss.n2824 dvss 0.00735484
R9288 dvss.n2821 dvss 0.00735484
R9289 dvss.n2820 dvss 0.00735484
R9290 dvss.n2819 dvss 0.00735484
R9291 dvss.n2816 dvss 0.00735484
R9292 dvss.n2815 dvss 0.00735484
R9293 dvss dvss.n1696 0.00735484
R9294 dvss.n2812 dvss 0.00735484
R9295 dvss.n2811 dvss 0.00735484
R9296 dvss.n2808 dvss 0.00735484
R9297 dvss.n2807 dvss 0.00735484
R9298 dvss dvss.n1702 0.00735484
R9299 dvss.n2803 dvss 0.00735484
R9300 dvss.n2802 dvss 0.00735484
R9301 dvss.n2799 dvss 0.00735484
R9302 dvss.n2795 dvss 0.00735484
R9303 dvss.n2794 dvss 0.00735484
R9304 dvss.n2791 dvss 0.00735484
R9305 dvss.n2790 dvss 0.00735484
R9306 dvss.n2789 dvss 0.00735484
R9307 dvss.n2785 dvss 0.00735484
R9308 dvss.n2784 dvss 0.00735484
R9309 dvss.n2781 dvss 0.00735484
R9310 dvss.n2780 dvss 0.00735484
R9311 dvss.n2779 dvss 0.00735484
R9312 dvss.n2776 dvss 0.00735484
R9313 dvss.n2775 dvss 0.00735484
R9314 dvss.n2774 dvss 0.00735484
R9315 dvss.n2771 dvss 0.00735484
R9316 dvss.n2770 dvss 0.00735484
R9317 dvss.n2769 dvss 0.00735484
R9318 dvss.n2766 dvss 0.00735484
R9319 dvss.n2765 dvss 0.00735484
R9320 dvss dvss.n1727 0.00735484
R9321 dvss.n2762 dvss 0.00735484
R9322 dvss.n2761 dvss 0.00735484
R9323 dvss.n2758 dvss 0.00735484
R9324 dvss.n2757 dvss 0.00735484
R9325 dvss dvss.n1733 0.00735484
R9326 dvss.n2753 dvss 0.00735484
R9327 dvss.n2752 dvss 0.00735484
R9328 dvss.n2749 dvss 0.00735484
R9329 dvss.n2745 dvss 0.00735484
R9330 dvss.n2744 dvss 0.00735484
R9331 dvss.n2741 dvss 0.00735484
R9332 dvss.n2740 dvss 0.00735484
R9333 dvss.n2739 dvss 0.00735484
R9334 dvss.n2735 dvss 0.00735484
R9335 dvss.n2734 dvss 0.00735484
R9336 dvss.n2731 dvss 0.00735484
R9337 dvss.n2730 dvss 0.00735484
R9338 dvss.n2729 dvss 0.00735484
R9339 dvss.n2726 dvss 0.00735484
R9340 dvss.n2725 dvss 0.00735484
R9341 dvss.n2724 dvss 0.00735484
R9342 dvss.n2721 dvss 0.00735484
R9343 dvss.n2720 dvss 0.00735484
R9344 dvss.n2719 dvss 0.00735484
R9345 dvss.n2716 dvss 0.00735484
R9346 dvss.n2715 dvss 0.00735484
R9347 dvss dvss.n1758 0.00735484
R9348 dvss.n2712 dvss 0.00735484
R9349 dvss.n2711 dvss 0.00735484
R9350 dvss.n2708 dvss 0.00735484
R9351 dvss.n2707 dvss 0.00735484
R9352 dvss dvss.n1764 0.00735484
R9353 dvss.n2703 dvss 0.00735484
R9354 dvss.n2702 dvss 0.00735484
R9355 dvss.n2699 dvss 0.00735484
R9356 dvss.n2695 dvss 0.00735484
R9357 dvss.n2694 dvss 0.00735484
R9358 dvss.n2691 dvss 0.00735484
R9359 dvss.n2690 dvss 0.00735484
R9360 dvss.n2689 dvss 0.00735484
R9361 dvss.n2685 dvss 0.00735484
R9362 dvss.n2684 dvss 0.00735484
R9363 dvss.n1775 dvss 0.00735484
R9364 dvss dvss.n3552 0.00735484
R9365 dvss dvss.n3553 0.00735484
R9366 dvss.n3567 dvss 0.00735484
R9367 dvss.n3566 dvss 0.00735484
R9368 dvss.n3565 dvss 0.00735484
R9369 dvss.n3562 dvss 0.00735484
R9370 dvss.n3561 dvss 0.00735484
R9371 dvss.n3560 dvss 0.00735484
R9372 dvss dvss.n3577 0.00735484
R9373 dvss dvss.n3578 0.00735484
R9374 dvss dvss.n3579 0.00735484
R9375 dvss.n3580 dvss 0.00735484
R9376 dvss.n3586 dvss 0.00735484
R9377 dvss.n3585 dvss 0.00735484
R9378 dvss.n3584 dvss 0.00735484
R9379 dvss dvss.n3594 0.00735484
R9380 dvss.n3596 dvss 0.00735484
R9381 dvss.n3595 dvss 0.00735484
R9382 dvss.n3601 dvss 0.00735484
R9383 dvss.n151 dvss 0.00735484
R9384 dvss dvss.n3609 0.00735484
R9385 dvss dvss.n3610 0.00735484
R9386 dvss.n3619 dvss 0.00735484
R9387 dvss.n3618 dvss 0.00735484
R9388 dvss.n3614 dvss 0.00735484
R9389 dvss dvss.n3627 0.00735484
R9390 dvss dvss.n3628 0.00735484
R9391 dvss.n3632 dvss 0.00735484
R9392 dvss.n3631 dvss 0.00735484
R9393 dvss.n3630 dvss 0.00735484
R9394 dvss.n3629 dvss 0.00735484
R9395 dvss dvss.n3643 0.00735484
R9396 dvss dvss.n783 0.00695161
R9397 dvss.n1159 dvss 0.00695161
R9398 dvss dvss.n1202 0.00695161
R9399 dvss.n1632 dvss 0.00695161
R9400 dvss dvss.n1675 0.00695161
R9401 dvss dvss.n1706 0.00695161
R9402 dvss dvss.n1737 0.00695161
R9403 dvss dvss.n1768 0.00695161
R9404 dvss dvss.n150 0.00695161
R9405 dvss dvss.n886 0.0064691
R9406 dvss.n888 dvss 0.0064691
R9407 dvss.n887 dvss 0.0064691
R9408 dvss dvss.n912 0.0064691
R9409 dvss dvss.n913 0.0064691
R9410 dvss.n919 dvss 0.0064691
R9411 dvss dvss.n929 0.0064691
R9412 dvss dvss.n930 0.0064691
R9413 dvss.n934 dvss 0.0064691
R9414 dvss.n937 dvss 0.0064691
R9415 dvss.n937 dvss 0.0064691
R9416 dvss.n936 dvss 0.0064691
R9417 dvss.n932 dvss 0.0064691
R9418 dvss.n931 dvss 0.0064691
R9419 dvss dvss.n949 0.0064691
R9420 dvss.n955 dvss 0.0064691
R9421 dvss.n954 dvss 0.0064691
R9422 dvss dvss.n963 0.0064691
R9423 dvss dvss.n964 0.0064691
R9424 dvss.n965 dvss 0.0064691
R9425 dvss.n973 dvss 0.0064691
R9426 dvss.n972 dvss 0.0064691
R9427 dvss.n978 dvss 0.0064691
R9428 dvss.n977 dvss 0.0064691
R9429 dvss.n755 dvss 0.0064691
R9430 dvss.n994 dvss 0.0064691
R9431 dvss.n993 dvss 0.0064691
R9432 dvss.n984 dvss 0.0064691
R9433 dvss.n738 dvss 0.0064691
R9434 dvss.n737 dvss 0.0064691
R9435 dvss.n1016 dvss 0.0064691
R9436 dvss.n1015 dvss 0.0064691
R9437 dvss.n1014 dvss 0.0064691
R9438 dvss.n1030 dvss 0.0064691
R9439 dvss.n1029 dvss 0.0064691
R9440 dvss.n1040 dvss 0.0064691
R9441 dvss.n1039 dvss 0.0064691
R9442 dvss dvss.n621 0.0064691
R9443 dvss dvss.n622 0.0064691
R9444 dvss dvss.n1049 0.0064691
R9445 dvss dvss.n1052 0.0064691
R9446 dvss.n1058 dvss 0.0064691
R9447 dvss.n1057 dvss 0.0064691
R9448 dvss dvss.n632 0.0064691
R9449 dvss.n709 dvss 0.0064691
R9450 dvss dvss.n633 0.0064691
R9451 dvss.n1068 dvss 0.0064691
R9452 dvss.n1067 dvss 0.0064691
R9453 dvss dvss.n640 0.0064691
R9454 dvss.n1071 dvss 0.0064691
R9455 dvss dvss.n641 0.0064691
R9456 dvss.n1075 dvss 0.0064691
R9457 dvss dvss.n642 0.0064691
R9458 dvss.n1080 dvss 0.0064691
R9459 dvss.n707 dvss 0.0064691
R9460 dvss dvss.n659 0.0064691
R9461 dvss.n704 dvss 0.0064691
R9462 dvss.n703 dvss 0.0064691
R9463 dvss.n702 dvss 0.0064691
R9464 dvss.n693 dvss 0.0064691
R9465 dvss.n690 dvss 0.0064691
R9466 dvss dvss.n1296 0.0064691
R9467 dvss.n1297 dvss 0.0064691
R9468 dvss dvss.n563 0.0064691
R9469 dvss.n1318 dvss 0.0064691
R9470 dvss.n1315 dvss 0.0064691
R9471 dvss.n1314 dvss 0.0064691
R9472 dvss dvss.n1328 0.0064691
R9473 dvss.n1329 dvss 0.0064691
R9474 dvss.n1334 dvss 0.0064691
R9475 dvss.n1342 dvss 0.0064691
R9476 dvss.n1341 dvss 0.0064691
R9477 dvss dvss.n1346 0.0064691
R9478 dvss.n1347 dvss 0.0064691
R9479 dvss dvss.n1354 0.0064691
R9480 dvss.n1355 dvss 0.0064691
R9481 dvss.n1362 dvss 0.0064691
R9482 dvss.n1361 dvss 0.0064691
R9483 dvss.n1366 dvss 0.0064691
R9484 dvss.n1365 dvss 0.0064691
R9485 dvss.n1383 dvss 0.0064691
R9486 dvss.n1382 dvss 0.0064691
R9487 dvss.n1393 dvss 0.0064691
R9488 dvss.n1392 dvss 0.0064691
R9489 dvss.n1391 dvss 0.0064691
R9490 dvss.n1407 dvss 0.0064691
R9491 dvss.n1406 dvss 0.0064691
R9492 dvss.n1416 dvss 0.0064691
R9493 dvss.n1415 dvss 0.0064691
R9494 dvss.n1574 dvss 0.0064691
R9495 dvss.n1573 dvss 0.0064691
R9496 dvss.n1572 dvss 0.0064691
R9497 dvss.n1569 dvss 0.0064691
R9498 dvss.n1568 dvss 0.0064691
R9499 dvss.n1567 dvss 0.0064691
R9500 dvss.n1564 dvss 0.0064691
R9501 dvss.n1436 dvss 0.0064691
R9502 dvss.n1561 dvss 0.0064691
R9503 dvss.n1560 dvss 0.0064691
R9504 dvss dvss.n1499 0.0064691
R9505 dvss.n1500 dvss 0.0064691
R9506 dvss.n1556 dvss 0.0064691
R9507 dvss.n1555 dvss 0.0064691
R9508 dvss.n1546 dvss 0.0064691
R9509 dvss.n1552 dvss 0.0064691
R9510 dvss.n1551 dvss 0.0064691
R9511 dvss.n1544 dvss 0.0064691
R9512 dvss dvss.n1457 0.0064691
R9513 dvss.n1541 dvss 0.0064691
R9514 dvss.n1540 dvss 0.0064691
R9515 dvss.n1539 dvss 0.0064691
R9516 dvss.n1530 dvss 0.0064691
R9517 dvss.n1527 dvss 0.0064691
R9518 dvss dvss.n2886 0.0064691
R9519 dvss.n2887 dvss 0.0064691
R9520 dvss.n2911 dvss 0.0064691
R9521 dvss.n2908 dvss 0.0064691
R9522 dvss.n2907 dvss 0.0064691
R9523 dvss.n2906 dvss 0.0064691
R9524 dvss dvss.n2920 0.0064691
R9525 dvss.n2921 dvss 0.0064691
R9526 dvss.n2926 dvss 0.0064691
R9527 dvss.n2934 dvss 0.0064691
R9528 dvss.n2933 dvss 0.0064691
R9529 dvss dvss.n2938 0.0064691
R9530 dvss.n2939 dvss 0.0064691
R9531 dvss dvss.n2946 0.0064691
R9532 dvss.n2947 dvss 0.0064691
R9533 dvss.n2954 dvss 0.0064691
R9534 dvss.n2953 dvss 0.0064691
R9535 dvss.n2958 dvss 0.0064691
R9536 dvss.n2957 dvss 0.0064691
R9537 dvss.n2975 dvss 0.0064691
R9538 dvss.n2974 dvss 0.0064691
R9539 dvss.n2985 dvss 0.0064691
R9540 dvss.n2984 dvss 0.0064691
R9541 dvss.n2983 dvss 0.0064691
R9542 dvss.n3000 dvss 0.0064691
R9543 dvss.n2999 dvss 0.0064691
R9544 dvss.n3009 dvss 0.0064691
R9545 dvss.n3008 dvss 0.0064691
R9546 dvss.n402 dvss 0.0064691
R9547 dvss.n3031 dvss 0.0064691
R9548 dvss.n3028 dvss 0.0064691
R9549 dvss.n3027 dvss 0.0064691
R9550 dvss dvss.n3039 0.0064691
R9551 dvss.n3040 dvss 0.0064691
R9552 dvss.n3048 dvss 0.0064691
R9553 dvss.n385 dvss 0.0064691
R9554 dvss.n384 dvss 0.0064691
R9555 dvss.n3060 dvss 0.0064691
R9556 dvss.n3059 dvss 0.0064691
R9557 dvss.n3071 dvss 0.0064691
R9558 dvss.n3070 dvss 0.0064691
R9559 dvss.n3074 dvss 0.0064691
R9560 dvss.n3066 dvss 0.0064691
R9561 dvss.n3065 dvss 0.0064691
R9562 dvss.n3083 dvss 0.0064691
R9563 dvss.n3091 dvss 0.0064691
R9564 dvss.n3090 dvss 0.0064691
R9565 dvss dvss.n3098 0.0064691
R9566 dvss.n3105 dvss 0.0064691
R9567 dvss.n3104 dvss 0.0064691
R9568 dvss.n3117 dvss 0.0064691
R9569 dvss.n3116 dvss 0.0064691
R9570 dvss.n3126 dvss 0.0064691
R9571 dvss.n3125 dvss 0.0064691
R9572 dvss.n3129 dvss 0.0064691
R9573 dvss.n3144 dvss 0.0064691
R9574 dvss.n3143 dvss 0.0064691
R9575 dvss.n3142 dvss 0.0064691
R9576 dvss dvss.n3153 0.0064691
R9577 dvss.n3154 dvss 0.0064691
R9578 dvss.n3165 dvss 0.0064691
R9579 dvss.n3164 dvss 0.0064691
R9580 dvss dvss.n3160 0.0064691
R9581 dvss.n3161 dvss 0.0064691
R9582 dvss.n3176 dvss 0.0064691
R9583 dvss dvss.n3179 0.0064691
R9584 dvss.n3180 dvss 0.0064691
R9585 dvss.n3187 dvss 0.0064691
R9586 dvss.n3186 dvss 0.0064691
R9587 dvss.n309 dvss 0.0064691
R9588 dvss.n3199 dvss 0.0064691
R9589 dvss.n3207 dvss 0.0064691
R9590 dvss.n3206 dvss 0.0064691
R9591 dvss dvss.n3214 0.0064691
R9592 dvss.n3221 dvss 0.0064691
R9593 dvss.n3220 dvss 0.0064691
R9594 dvss.n3233 dvss 0.0064691
R9595 dvss.n3232 dvss 0.0064691
R9596 dvss.n3242 dvss 0.0064691
R9597 dvss.n3241 dvss 0.0064691
R9598 dvss.n3245 dvss 0.0064691
R9599 dvss.n3260 dvss 0.0064691
R9600 dvss.n3259 dvss 0.0064691
R9601 dvss.n3258 dvss 0.0064691
R9602 dvss dvss.n3268 0.0064691
R9603 dvss.n3269 dvss 0.0064691
R9604 dvss.n3283 dvss 0.0064691
R9605 dvss.n3282 dvss 0.0064691
R9606 dvss dvss.n3278 0.0064691
R9607 dvss.n3279 dvss 0.0064691
R9608 dvss dvss.n3293 0.0064691
R9609 dvss dvss.n3294 0.0064691
R9610 dvss.n3295 dvss 0.0064691
R9611 dvss.n3306 dvss 0.0064691
R9612 dvss dvss.n3301 0.0064691
R9613 dvss.n3303 dvss 0.0064691
R9614 dvss.n3302 dvss 0.0064691
R9615 dvss.n3323 dvss 0.0064691
R9616 dvss.n3322 dvss 0.0064691
R9617 dvss.n3333 dvss 0.0064691
R9618 dvss.n3332 dvss 0.0064691
R9619 dvss.n3331 dvss 0.0064691
R9620 dvss.n3347 dvss 0.0064691
R9621 dvss.n3346 dvss 0.0064691
R9622 dvss.n3356 dvss 0.0064691
R9623 dvss.n3355 dvss 0.0064691
R9624 dvss.n3540 dvss 0.0064691
R9625 dvss.n3539 dvss 0.0064691
R9626 dvss.n3538 dvss 0.0064691
R9627 dvss.n3535 dvss 0.0064691
R9628 dvss.n3534 dvss 0.0064691
R9629 dvss.n3533 dvss 0.0064691
R9630 dvss.n3530 dvss 0.0064691
R9631 dvss.n3376 dvss 0.0064691
R9632 dvss.n3527 dvss 0.0064691
R9633 dvss.n3526 dvss 0.0064691
R9634 dvss dvss.n3426 0.0064691
R9635 dvss.n3427 dvss 0.0064691
R9636 dvss.n3522 dvss 0.0064691
R9637 dvss.n3521 dvss 0.0064691
R9638 dvss.n3512 dvss 0.0064691
R9639 dvss.n3518 dvss 0.0064691
R9640 dvss.n3517 dvss 0.0064691
R9641 dvss.n3510 dvss 0.0064691
R9642 dvss.n3401 dvss 0.0064691
R9643 dvss.n3507 dvss 0.0064691
R9644 dvss.n3506 dvss 0.0064691
R9645 dvss.n3505 dvss 0.0064691
R9646 dvss.n3475 dvss 0.0064691
R9647 dvss.n3418 dvss 0.0064691
R9648 dvss.n3417 dvss 0.0064691
R9649 dvss dvss.n3404 0.0064691
R9650 dvss.n3491 dvss 0.0064691
R9651 dvss.n3490 dvss 0.0064691
R9652 dvss.n3646 dvss 0.0064691
R9653 dvss.n2625 dvss.n2000 0.00641216
R9654 dvss.n2578 dvss.n2033 0.00641216
R9655 dvss.n2531 dvss.n2069 0.00641216
R9656 dvss.n2484 dvss.n2105 0.00641216
R9657 dvss.n2437 dvss.n2141 0.00641216
R9658 dvss.n2390 dvss.n2177 0.00641216
R9659 dvss.n2343 dvss.n2209 0.00641216
R9660 dvss.n2296 dvss.n2295 0.00641216
R9661 dvss.n3694 dvss.n95 0.00641216
R9662 dvss.n913 dvss 0.00611798
R9663 dvss.n1000 dvss 0.00611798
R9664 dvss dvss.n651 0.00611798
R9665 dvss.n1378 dvss 0.00611798
R9666 dvss dvss.n1448 0.00611798
R9667 dvss.n2970 dvss 0.00611798
R9668 dvss.n3086 dvss 0.00611798
R9669 dvss.n3202 dvss 0.00611798
R9670 dvss.n3318 dvss 0.00611798
R9671 dvss dvss.n3388 0.00611798
R9672 dvss.n918 dvss.n917 0.00576685
R9673 dvss.n811 dvss 0.00574194
R9674 dvss.n1170 dvss 0.00574194
R9675 dvss dvss.n1249 0.00574194
R9676 dvss.n1643 dvss 0.00574194
R9677 dvss dvss.n2839 0.00574194
R9678 dvss dvss.n2789 0.00574194
R9679 dvss dvss.n2739 0.00574194
R9680 dvss dvss.n2689 0.00574194
R9681 dvss dvss.n3618 0.00574194
R9682 dvss dvss.n2646 0.00556757
R9683 dvss dvss.n954 0.00541573
R9684 dvss.n998 dvss 0.00541573
R9685 dvss dvss.n1057 0.00541573
R9686 dvss.n708 dvss 0.00541573
R9687 dvss.n1329 dvss 0.00541573
R9688 dvss dvss.n1381 0.00541573
R9689 dvss dvss.n1567 0.00541573
R9690 dvss.n1545 dvss 0.00541573
R9691 dvss.n2921 dvss 0.00541573
R9692 dvss dvss.n2973 0.00541573
R9693 dvss.n3040 dvss 0.00541573
R9694 dvss dvss.n3089 0.00541573
R9695 dvss.n3154 dvss 0.00541573
R9696 dvss dvss.n3205 0.00541573
R9697 dvss.n3269 dvss 0.00541573
R9698 dvss dvss.n3321 0.00541573
R9699 dvss dvss.n3533 0.00541573
R9700 dvss.n3511 dvss 0.00541573
R9701 dvss dvss.n1014 0.00506461
R9702 dvss dvss.n620 0.00506461
R9703 dvss dvss.n702 0.00506461
R9704 dvss.n1300 dvss 0.00506461
R9705 dvss dvss.n1391 0.00506461
R9706 dvss.n1577 dvss 0.00506461
R9707 dvss dvss.n1539 0.00506461
R9708 dvss.n2890 dvss 0.00506461
R9709 dvss dvss.n2983 0.00506461
R9710 dvss.n3012 dvss 0.00506461
R9711 dvss dvss.n3104 0.00506461
R9712 dvss.n3130 dvss 0.00506461
R9713 dvss dvss.n3220 0.00506461
R9714 dvss.n3246 dvss 0.00506461
R9715 dvss dvss.n3331 0.00506461
R9716 dvss.n3543 dvss 0.00506461
R9717 dvss dvss.n3505 0.00506461
R9718 dvss.n3494 dvss 0.00506461
R9719 dvss.n813 dvss 0.00493548
R9720 dvss.n1173 dvss 0.00493548
R9721 dvss.n1246 dvss 0.00493548
R9722 dvss.n1646 dvss 0.00493548
R9723 dvss.n2836 dvss 0.00493548
R9724 dvss.n2786 dvss 0.00493548
R9725 dvss.n2736 dvss 0.00493548
R9726 dvss.n2686 dvss 0.00493548
R9727 dvss.n3615 dvss 0.00493548
R9728 dvss.n952 dvss 0.00401124
R9729 dvss.n1009 dvss.n722 0.00401124
R9730 dvss.n1055 dvss 0.00401124
R9731 dvss.n698 dvss.n694 0.00401124
R9732 dvss dvss.n1333 0.00401124
R9733 dvss.n1386 dvss.n516 0.00401124
R9734 dvss.n1565 dvss 0.00401124
R9735 dvss.n1535 dvss.n1531 0.00401124
R9736 dvss dvss.n2925 0.00401124
R9737 dvss.n2978 dvss.n407 0.00401124
R9738 dvss.n3044 dvss 0.00401124
R9739 dvss.n3099 dvss.n344 0.00401124
R9740 dvss dvss.n3158 0.00401124
R9741 dvss.n3215 dvss.n280 0.00401124
R9742 dvss.n3273 dvss 0.00401124
R9743 dvss.n3326 dvss.n217 0.00401124
R9744 dvss.n3531 dvss 0.00401124
R9745 dvss.n3501 dvss.n3400 0.00401124
R9746 dvss.n2658 dvss 0.00387838
R9747 dvss.n2602 dvss.n2019 0.00387838
R9748 dvss.n2591 dvss.n2590 0.00387838
R9749 dvss.n2555 dvss.n2055 0.00387838
R9750 dvss.n2544 dvss.n2543 0.00387838
R9751 dvss.n2508 dvss.n2091 0.00387838
R9752 dvss.n2497 dvss.n2496 0.00387838
R9753 dvss.n2461 dvss.n2127 0.00387838
R9754 dvss.n2450 dvss.n2449 0.00387838
R9755 dvss.n2414 dvss.n2163 0.00387838
R9756 dvss.n2403 dvss.n2402 0.00387838
R9757 dvss.n2367 dvss.n2197 0.00387838
R9758 dvss.n2356 dvss.n2355 0.00387838
R9759 dvss.n2320 dvss.n2252 0.00387838
R9760 dvss.n2309 dvss.n2308 0.00387838
R9761 dvss.n3718 dvss.n83 0.00387838
R9762 dvss.n3707 dvss.n3706 0.00387838
R9763 dvss.n3671 dvss.n111 0.00387838
R9764 dvss.n3660 dvss.n3659 0.00387838
R9765 dvss dvss.n778 0.00372581
R9766 dvss.n803 dvss 0.00372581
R9767 dvss dvss.n599 0.00372581
R9768 dvss dvss.n590 0.00372581
R9769 dvss.n1198 dvss 0.00372581
R9770 dvss dvss.n1254 0.00372581
R9771 dvss dvss.n489 0.00372581
R9772 dvss dvss.n480 0.00372581
R9773 dvss.n1671 dvss 0.00372581
R9774 dvss dvss.n2844 0.00372581
R9775 dvss.n1702 dvss 0.00372581
R9776 dvss dvss.n2794 0.00372581
R9777 dvss.n1733 dvss 0.00372581
R9778 dvss dvss.n2744 0.00372581
R9779 dvss.n1764 dvss 0.00372581
R9780 dvss dvss.n2694 0.00372581
R9781 dvss.n3594 dvss 0.00372581
R9782 dvss.n3609 dvss 0.00372581
R9783 dvss.n910 dvss.n909 0.00366011
R9784 dvss.n928 dvss.n868 0.00366011
R9785 dvss.n909 dvss 0.00330899
R9786 dvss dvss.n928 0.00330899
R9787 dvss dvss.n755 0.00330899
R9788 dvss dvss.n738 0.00330899
R9789 dvss dvss.n641 0.00330899
R9790 dvss dvss.n707 0.00330899
R9791 dvss.n1362 dvss 0.00330899
R9792 dvss.n1383 dvss 0.00330899
R9793 dvss dvss.n1555 0.00330899
R9794 dvss dvss.n1544 0.00330899
R9795 dvss.n2954 dvss 0.00330899
R9796 dvss.n2975 dvss 0.00330899
R9797 dvss.n3074 dvss 0.00330899
R9798 dvss.n3091 dvss 0.00330899
R9799 dvss.n3187 dvss 0.00330899
R9800 dvss.n3207 dvss 0.00330899
R9801 dvss.n3306 dvss 0.00330899
R9802 dvss.n3323 dvss 0.00330899
R9803 dvss dvss.n3521 0.00330899
R9804 dvss dvss.n3510 0.00330899
R9805 dvss dvss.n2593 0.00303378
R9806 dvss dvss.n2546 0.00303378
R9807 dvss dvss.n2499 0.00303378
R9808 dvss dvss.n2452 0.00303378
R9809 dvss dvss.n2405 0.00303378
R9810 dvss dvss.n2358 0.00303378
R9811 dvss dvss.n2311 0.00303378
R9812 dvss dvss.n3709 0.00303378
R9813 dvss dvss.n3662 0.00303378
R9814 dvss.n952 dvss.n763 0.00295787
R9815 dvss.n725 dvss 0.00295787
R9816 dvss.n1009 dvss 0.00295787
R9817 dvss.n1055 dvss.n631 0.00295787
R9818 dvss.n699 dvss 0.00295787
R9819 dvss.n694 dvss 0.00295787
R9820 dvss.n1333 dvss.n552 0.00295787
R9821 dvss.n519 dvss 0.00295787
R9822 dvss.n1386 dvss 0.00295787
R9823 dvss.n1565 dvss.n1429 0.00295787
R9824 dvss.n1536 dvss 0.00295787
R9825 dvss.n1531 dvss 0.00295787
R9826 dvss.n2925 dvss.n443 0.00295787
R9827 dvss.n410 dvss 0.00295787
R9828 dvss.n2978 dvss 0.00295787
R9829 dvss.n3045 dvss.n3044 0.00295787
R9830 dvss.n347 dvss 0.00295787
R9831 dvss.n3099 dvss 0.00295787
R9832 dvss.n3158 dvss.n319 0.00295787
R9833 dvss.n283 dvss 0.00295787
R9834 dvss.n3215 dvss 0.00295787
R9835 dvss.n3274 dvss.n3273 0.00295787
R9836 dvss.n220 dvss 0.00295787
R9837 dvss.n3326 dvss 0.00295787
R9838 dvss.n3531 dvss.n3369 0.00295787
R9839 dvss.n3502 dvss 0.00295787
R9840 dvss dvss.n3400 0.00295787
R9841 dvss.n789 dvss 0.00291935
R9842 dvss.n813 dvss.n810 0.00291935
R9843 dvss.n1139 dvss 0.00291935
R9844 dvss.n1174 dvss.n1173 0.00291935
R9845 dvss.n1272 dvss 0.00291935
R9846 dvss.n1246 dvss.n1208 0.00291935
R9847 dvss.n1612 dvss 0.00291935
R9848 dvss.n1647 dvss.n1646 0.00291935
R9849 dvss.n2862 dvss 0.00291935
R9850 dvss.n2836 dvss.n1681 0.00291935
R9851 dvss.n2812 dvss 0.00291935
R9852 dvss.n2786 dvss.n1712 0.00291935
R9853 dvss.n2762 dvss 0.00291935
R9854 dvss.n2736 dvss.n1743 0.00291935
R9855 dvss.n2712 dvss 0.00291935
R9856 dvss.n2686 dvss.n1774 0.00291935
R9857 dvss.n3580 dvss 0.00291935
R9858 dvss.n3615 dvss.n3613 0.00291935
R9859 dvss.n973 dvss 0.00260674
R9860 dvss.n1033 dvss.n725 0.00260674
R9861 dvss.n1068 dvss 0.00260674
R9862 dvss.n699 dvss.n664 0.00260674
R9863 dvss.n1346 dvss 0.00260674
R9864 dvss.n1410 dvss.n519 0.00260674
R9865 dvss dvss.n1560 0.00260674
R9866 dvss.n1536 dvss.n1462 0.00260674
R9867 dvss.n2938 dvss 0.00260674
R9868 dvss.n3003 dvss.n410 0.00260674
R9869 dvss.n3060 dvss 0.00260674
R9870 dvss.n3120 dvss.n347 0.00260674
R9871 dvss.n3161 dvss 0.00260674
R9872 dvss.n3236 dvss.n283 0.00260674
R9873 dvss.n3279 dvss 0.00260674
R9874 dvss.n3350 dvss.n220 0.00260674
R9875 dvss dvss.n3526 0.00260674
R9876 dvss.n3502 dvss.n3399 0.00260674
R9877 dvss dvss.n885 0.00190449
R9878 dvss.n1034 dvss.n1033 0.00190449
R9879 dvss.n1037 dvss.n620 0.00190449
R9880 dvss.n696 dvss.n664 0.00190449
R9881 dvss.n1300 dvss.n1299 0.00190449
R9882 dvss.n1411 dvss.n1410 0.00190449
R9883 dvss.n1577 dvss.n511 0.00190449
R9884 dvss.n1533 dvss.n1462 0.00190449
R9885 dvss.n2890 dvss.n2889 0.00190449
R9886 dvss.n3004 dvss.n3003 0.00190449
R9887 dvss.n3012 dvss.n401 0.00190449
R9888 dvss.n3121 dvss.n3120 0.00190449
R9889 dvss.n3130 dvss.n339 0.00190449
R9890 dvss.n3237 dvss.n3236 0.00190449
R9891 dvss.n3246 dvss.n275 0.00190449
R9892 dvss.n3351 dvss.n3350 0.00190449
R9893 dvss.n3543 dvss.n212 0.00190449
R9894 dvss.n3499 dvss.n3399 0.00190449
R9895 dvss.n3495 dvss.n3494 0.00190449
R9896 dvss.n999 dvss.n998 0.00155337
R9897 dvss dvss.n1039 0.00155337
R9898 dvss.n708 dvss.n652 0.00155337
R9899 dvss.n1297 dvss 0.00155337
R9900 dvss.n1381 dvss.n532 0.00155337
R9901 dvss dvss.n1415 0.00155337
R9902 dvss.n1545 dvss.n1449 0.00155337
R9903 dvss.n2887 dvss 0.00155337
R9904 dvss.n2973 dvss.n423 0.00155337
R9905 dvss dvss.n3008 0.00155337
R9906 dvss.n3089 dvss.n363 0.00155337
R9907 dvss dvss.n3125 0.00155337
R9908 dvss.n3205 dvss.n299 0.00155337
R9909 dvss dvss.n3241 0.00155337
R9910 dvss.n3321 dvss.n233 0.00155337
R9911 dvss dvss.n3355 0.00155337
R9912 dvss.n3511 dvss.n3389 0.00155337
R9913 dvss dvss.n3404 0.00155337
R9914 dvss.n2644 dvss.n2643 0.00134459
R9915 dvss.n917 dvss 0.00120225
R9916 dvss.n800 dvss.n783 0.000903226
R9917 dvss.n818 dvss 0.000903226
R9918 dvss.n1159 dvss.n589 0.000903226
R9919 dvss dvss.n582 0.000903226
R9920 dvss.n1258 dvss.n1202 0.000903226
R9921 dvss dvss.n1244 0.000903226
R9922 dvss.n1632 dvss.n479 0.000903226
R9923 dvss dvss.n472 0.000903226
R9924 dvss.n2848 dvss.n1675 0.000903226
R9925 dvss dvss.n2834 0.000903226
R9926 dvss.n2798 dvss.n1706 0.000903226
R9927 dvss dvss.n2784 0.000903226
R9928 dvss.n2748 dvss.n1737 0.000903226
R9929 dvss dvss.n2734 0.000903226
R9930 dvss.n2698 dvss.n1768 0.000903226
R9931 dvss dvss.n2684 0.000903226
R9932 dvss.n3600 dvss.n150 0.000903226
R9933 dvss.n3627 dvss 0.000903226
R9934 dvss.n1000 dvss.n742 0.000851124
R9935 dvss.n1030 dvss 0.000851124
R9936 dvss.n1079 dvss.n651 0.000851124
R9937 dvss dvss.n693 0.000851124
R9938 dvss.n1379 dvss.n1378 0.000851124
R9939 dvss.n1407 dvss 0.000851124
R9940 dvss.n1550 dvss.n1448 0.000851124
R9941 dvss dvss.n1530 0.000851124
R9942 dvss.n2971 dvss.n2970 0.000851124
R9943 dvss.n3000 dvss 0.000851124
R9944 dvss.n3087 dvss.n3086 0.000851124
R9945 dvss.n3117 dvss 0.000851124
R9946 dvss.n3203 dvss.n3202 0.000851124
R9947 dvss.n3233 dvss 0.000851124
R9948 dvss.n3319 dvss.n3318 0.000851124
R9949 dvss.n3347 dvss 0.000851124
R9950 dvss.n3516 dvss.n3388 0.000851124
R9951 dvss.n3475 dvss 0.000851124
R9952 avdd.n1200 avdd.n1199 113249
R9953 avdd.n1199 avdd.n1198 85895.3
R9954 avdd.n1200 avdd.n1167 82364.3
R9955 avdd.n1201 avdd.n1166 55683.2
R9956 avdd.n1198 avdd.n1168 54827.6
R9957 avdd.n1181 avdd.n1167 54152.8
R9958 avdd.n1182 avdd.n1168 47563.1
R9959 avdd.n1197 avdd.n1166 42329.2
R9960 avdd.n1201 avdd.n1165 40605.4
R9961 avdd.n1197 avdd.n1169 27162.2
R9962 avdd.n1179 avdd.n1165 26862.2
R9963 avdd.n1180 avdd.n1169 23168.1
R9964 avdd.n1183 avdd.n1181 23082.1
R9965 avdd.n1081 avdd.n1080 22451.2
R9966 avdd.n1082 avdd.n1081 22451.2
R9967 avdd.n1082 avdd.n1078 22451.2
R9968 avdd.n1080 avdd.n1078 22451.2
R9969 avdd.n1183 avdd.n1182 16349.3
R9970 avdd.n1230 avdd.n1223 13391.1
R9971 avdd.n1230 avdd.n1224 13391.1
R9972 avdd.n1265 avdd.n1224 13391.1
R9973 avdd.n1265 avdd.n1223 13391.1
R9974 avdd.n1146 avdd.n951 12351.3
R9975 avdd.n975 avdd.n951 12351.3
R9976 avdd.n1184 avdd.n1179 11693.5
R9977 avdd.n1079 avdd.n1077 11356.2
R9978 avdd.n1083 avdd.n1077 11356.2
R9979 avdd.n1083 avdd.n1076 11356.2
R9980 avdd.n1079 avdd.n1076 11356.2
R9981 avdd.n1142 avdd.n954 10507.7
R9982 avdd.n1142 avdd.n950 10507.7
R9983 avdd.n1144 avdd.n952 10039.9
R9984 avdd.n1145 avdd.n1144 10039.9
R9985 avdd.n1196 avdd.n1171 9834.54
R9986 avdd.n1350 avdd.n679 9739.14
R9987 avdd.n1350 avdd.n680 9739.14
R9988 avdd.n1349 avdd.n680 9739.14
R9989 avdd.n1349 avdd.n679 9739.14
R9990 avdd.n1192 avdd.n1171 8773.65
R9991 avdd.n1184 avdd.n1180 7929.73
R9992 avdd.n1196 avdd.n1170 6313.41
R9993 avdd.n1177 avdd.n1176 6233.98
R9994 avdd.n1189 avdd.n1188 5357.93
R9995 avdd.n1174 avdd.n1163 4394.54
R9996 avdd.n1334 avdd.n1333 4316.28
R9997 avdd.n1336 avdd.n1333 4316.28
R9998 avdd.n1334 avdd.n1330 4316.28
R9999 avdd.n1336 avdd.n1330 4316.28
R10000 avdd.n1204 avdd.n1203 3955.2
R10001 avdd.n1301 avdd.n1216 3160.55
R10002 avdd.n1302 avdd.n1216 3160.55
R10003 avdd.n1202 avdd.n1164 3056.94
R10004 avdd.n1185 avdd.n1178 2722.26
R10005 avdd.n1084 avdd.n965 2632.66
R10006 avdd.n1075 avdd.n964 2621.36
R10007 avdd.n1264 avdd.n1225 2567.82
R10008 avdd.n1231 avdd.n1225 2567.82
R10009 avdd.n1085 avdd.n1074 2564.89
R10010 avdd.n1135 avdd.n1134 2540.05
R10011 avdd.n1232 avdd.n1226 2537.41
R10012 avdd.n1263 avdd.n1226 2537.41
R10013 avdd.n1295 avdd.n1267 2513.9
R10014 avdd.n1295 avdd.n1215 2513.9
R10015 avdd.n1296 avdd.n1220 2513.9
R10016 avdd.n1296 avdd.n1217 2513.9
R10017 avdd.n990 avdd.n973 2480.48
R10018 avdd.n988 avdd.n973 2480.48
R10019 avdd.n990 avdd.n974 2480.48
R10020 avdd.n988 avdd.n974 2480.48
R10021 avdd.n1290 avdd.n1284 2346.83
R10022 avdd.n1289 avdd.n1284 2346.83
R10023 avdd.n1019 avdd.n968 2342.02
R10024 avdd.n1146 avdd.n1145 2311.45
R10025 avdd.n975 avdd.n952 2311.45
R10026 avdd.n1015 avdd.n949 2059.86
R10027 avdd.n1149 avdd.n949 2059.86
R10028 avdd.n1149 avdd.n948 2059.86
R10029 avdd.n1015 avdd.n948 2059.86
R10030 avdd.n1141 avdd.n956 2000.19
R10031 avdd.n1141 avdd.n955 2000.19
R10032 avdd.n1019 avdd.n1018 1894.78
R10033 avdd.n1185 avdd.n1172 1848.47
R10034 avdd.n1302 avdd.n1215 1837.76
R10035 avdd.n1301 avdd.n1217 1837.76
R10036 avdd.n681 avdd.n677 1616.56
R10037 avdd.n1347 avdd.n682 1616.56
R10038 avdd.n682 avdd.n678 1616.56
R10039 avdd.n1352 avdd.n677 1615.06
R10040 avdd.n1286 avdd.n1220 1322.79
R10041 avdd.n1286 avdd.n1267 1322.79
R10042 avdd.n1221 avdd.n1217 1322.79
R10043 avdd.n1221 avdd.n1215 1322.79
R10044 avdd.n1064 avdd.n953 1237.08
R10045 avdd.n1126 avdd.n953 1237.08
R10046 avdd.n1192 avdd.n1164 1027.39
R10047 avdd.n1290 avdd.n1267 1024.03
R10048 avdd.n1289 avdd.n1220 1024.03
R10049 avdd.n1203 avdd.n1202 897.883
R10050 avdd.n1338 avdd.n1337 831.247
R10051 avdd.n1338 avdd.n1329 831.247
R10052 avdd.n73 avdd.t298 692.692
R10053 avdd avdd.t297 688.231
R10054 avdd.n1332 avdd.n1331 682.918
R10055 avdd.n1332 avdd.n1312 682.918
R10056 avdd.n1057 avdd.t110 660.24
R10057 avdd.t161 avdd.n1052 660.24
R10058 avdd.t85 avdd.n1049 660.24
R10059 avdd.n1046 avdd.t145 660.24
R10060 avdd.n1043 avdd.t169 660.24
R10061 avdd.t94 avdd.n1038 660.24
R10062 avdd.t117 avdd.n1035 660.24
R10063 avdd.n1032 avdd.t174 660.24
R10064 avdd.t105 avdd.n1027 660.24
R10065 avdd.n940 avdd.t135 660.24
R10066 avdd.n1106 avdd.t88 660.24
R10067 avdd.n1108 avdd.t115 660.24
R10068 avdd.n1110 avdd.t172 660.24
R10069 avdd.n1112 avdd.t97 660.24
R10070 avdd.n1114 avdd.t120 660.24
R10071 avdd.n1116 avdd.t148 660.24
R10072 avdd.n1118 avdd.t108 660.24
R10073 avdd.n1120 avdd.t130 660.24
R10074 avdd.n335 avdd.t382 648.668
R10075 avdd.n307 avdd.t326 648.668
R10076 avdd.n279 avdd.t352 648.668
R10077 avdd.n251 avdd.t374 648.668
R10078 avdd.n223 avdd.t273 648.668
R10079 avdd.n195 avdd.t317 648.668
R10080 avdd.n167 avdd.t287 648.668
R10081 avdd.n139 avdd.t378 648.668
R10082 avdd.n111 avdd.t359 648.668
R10083 avdd.n657 avdd.t314 648.668
R10084 avdd.n629 avdd.t7 648.668
R10085 avdd.n601 avdd.t1 648.668
R10086 avdd.n573 avdd.t75 648.668
R10087 avdd.n545 avdd.t196 648.668
R10088 avdd.n517 avdd.t291 648.668
R10089 avdd.n489 avdd.t259 648.668
R10090 avdd.n461 avdd.t252 648.668
R10091 avdd.n433 avdd.t241 648.668
R10092 avdd.n909 avdd.n692 624.808
R10093 avdd.n907 avdd.n693 624.808
R10094 avdd.n896 avdd.n895 624.808
R10095 avdd.n884 avdd.n712 624.808
R10096 avdd.n882 avdd.n713 624.808
R10097 avdd.n871 avdd.n870 624.808
R10098 avdd.n859 avdd.n732 624.808
R10099 avdd.n857 avdd.n733 624.808
R10100 avdd.n846 avdd.n845 624.808
R10101 avdd.n834 avdd.n752 624.808
R10102 avdd.n832 avdd.n753 624.808
R10103 avdd.n821 avdd.n820 624.808
R10104 avdd.n809 avdd.n772 624.808
R10105 avdd.n807 avdd.n773 624.808
R10106 avdd.n796 avdd.n795 624.808
R10107 avdd.n1065 avdd.n1064 612.894
R10108 avdd.n1126 avdd.n1125 612.894
R10109 avdd.n1300 avdd.n1213 609.883
R10110 avdd.n1014 avdd.n1013 598.801
R10111 avdd.n1012 avdd.n1011 598.801
R10112 avdd.n1010 avdd.n1009 598.801
R10113 avdd.n1008 avdd.n1007 598.801
R10114 avdd.n1006 avdd.n1005 598.801
R10115 avdd.n1004 avdd.n1003 598.801
R10116 avdd.n1002 avdd.n1001 598.801
R10117 avdd.n1000 avdd.n999 598.801
R10118 avdd.n998 avdd.n997 598.801
R10119 avdd.n1089 avdd.n1088 598.801
R10120 avdd.n1091 avdd.n1090 598.801
R10121 avdd.n1093 avdd.n1092 598.801
R10122 avdd.n1095 avdd.n1094 598.801
R10123 avdd.n1097 avdd.n1096 598.801
R10124 avdd.n1099 avdd.n1098 598.801
R10125 avdd.n1101 avdd.n1100 598.801
R10126 avdd.n1103 avdd.n1102 598.801
R10127 avdd.n1105 avdd.n1104 598.801
R10128 avdd.n1056 avdd.n1055 598.801
R10129 avdd.n1054 avdd.n1053 598.801
R10130 avdd.n1051 avdd.n1050 598.801
R10131 avdd.n1045 avdd.n1025 598.801
R10132 avdd.n1042 avdd.n1041 598.801
R10133 avdd.n1040 avdd.n1039 598.801
R10134 avdd.n1037 avdd.n1036 598.801
R10135 avdd.n1031 avdd.n1030 598.801
R10136 avdd.n1029 avdd.n1028 598.801
R10137 avdd.n1304 avdd.n1303 555.672
R10138 avdd.t46 avdd.t44 511.356
R10139 avdd.t50 avdd.t46 511.356
R10140 avdd.t362 avdd.t137 511.356
R10141 avdd.t364 avdd.t362 511.356
R10142 avdd.t154 avdd.t364 511.356
R10143 avdd.t366 avdd.t154 511.356
R10144 avdd.t368 avdd.t366 511.356
R10145 avdd.t99 avdd.t368 511.356
R10146 avdd.t84 avdd.t12 502.586
R10147 avdd.t12 avdd.t14 502.586
R10148 avdd.t21 avdd.t17 502.586
R10149 avdd.t17 avdd.t80 502.586
R10150 avdd.n667 avdd.t332 499.882
R10151 avdd.t344 avdd.t342 484.288
R10152 avdd.t213 avdd.t340 484.288
R10153 avdd.n1294 avdd.n1292 481.507
R10154 avdd.n1297 avdd.n1219 481.507
R10155 avdd.n987 avdd.n972 479.625
R10156 avdd.n991 avdd.n972 479.625
R10157 avdd.t44 avdd.t48 475.098
R10158 avdd.n954 avdd.n952 467.793
R10159 avdd.n1145 avdd.n950 467.793
R10160 avdd.n1288 avdd.n1283 454.024
R10161 avdd.n1018 avdd.n944 447.248
R10162 avdd.n1149 avdd.t213 437.699
R10163 avdd.n992 avdd.n971 437.082
R10164 avdd.n986 avdd.n971 437.082
R10165 avdd.n1291 avdd.n1283 423.818
R10166 avdd.n1016 avdd.n947 399.06
R10167 avdd.n1150 avdd.n947 399.06
R10168 avdd.n1271 avdd.t141 397.264
R10169 avdd.n1272 avdd.t149 397.135
R10170 avdd.n1273 avdd.t77 397.135
R10171 avdd.n676 avdd.t91 388.149
R10172 avdd.n920 avdd.t151 388.149
R10173 avdd.n921 avdd.t179 388.149
R10174 avdd.n922 avdd.t175 388.149
R10175 avdd.n923 avdd.t124 388.149
R10176 avdd.n924 avdd.t164 388.149
R10177 avdd.n925 avdd.t156 388.149
R10178 avdd.n926 avdd.t166 388.149
R10179 avdd.n928 avdd.t177 388.149
R10180 avdd.n929 avdd.t102 388.149
R10181 avdd.n930 avdd.t162 388.149
R10182 avdd.n931 avdd.t111 388.149
R10183 avdd.n932 avdd.t139 388.149
R10184 avdd.n933 avdd.t89 388.149
R10185 avdd.n934 avdd.t126 388.149
R10186 avdd.n331 avdd.t329 372.885
R10187 avdd.n303 avdd.t190 372.885
R10188 avdd.n275 avdd.t11 372.885
R10189 avdd.n247 avdd.t331 372.885
R10190 avdd.n219 avdd.t283 372.885
R10191 avdd.n191 avdd.t254 372.885
R10192 avdd.n163 avdd.t249 372.885
R10193 avdd.n135 avdd.t304 372.885
R10194 avdd.n107 avdd.t261 372.885
R10195 avdd.n653 avdd.t277 372.885
R10196 avdd.n625 avdd.t192 372.885
R10197 avdd.n597 avdd.t306 372.885
R10198 avdd.n569 avdd.t295 372.885
R10199 avdd.n541 avdd.t184 372.885
R10200 avdd.n513 avdd.t371 372.885
R10201 avdd.n485 avdd.t293 372.885
R10202 avdd.n457 avdd.t308 372.885
R10203 avdd.n429 avdd.t256 372.885
R10204 avdd.n1063 avdd.n1062 359.529
R10205 avdd.t185 avdd.n684 354.904
R10206 avdd.n1303 avdd.n1214 352
R10207 avdd.n1300 avdd.n1299 352
R10208 avdd.n1230 avdd.t99 345.817
R10209 avdd.n1015 avdd.t344 343.495
R10210 avdd.n1293 avdd.n1214 325.647
R10211 avdd.n1299 avdd.n1298 325.647
R10212 avdd.n990 avdd.t52 323.445
R10213 avdd.t246 avdd.n988 323.445
R10214 avdd.n324 avdd.n6 321.882
R10215 avdd.n310 avdd.n309 321.882
R10216 avdd.n4 avdd.n2 321.882
R10217 avdd.n296 avdd.n14 321.882
R10218 avdd.n282 avdd.n281 321.882
R10219 avdd.n12 avdd.n10 321.882
R10220 avdd.n268 avdd.n22 321.882
R10221 avdd.n254 avdd.n253 321.882
R10222 avdd.n20 avdd.n18 321.882
R10223 avdd.n240 avdd.n30 321.882
R10224 avdd.n226 avdd.n225 321.882
R10225 avdd.n28 avdd.n26 321.882
R10226 avdd.n212 avdd.n38 321.882
R10227 avdd.n198 avdd.n197 321.882
R10228 avdd.n36 avdd.n34 321.882
R10229 avdd.n184 avdd.n46 321.882
R10230 avdd.n170 avdd.n169 321.882
R10231 avdd.n44 avdd.n42 321.882
R10232 avdd.n156 avdd.n54 321.882
R10233 avdd.n142 avdd.n141 321.882
R10234 avdd.n52 avdd.n50 321.882
R10235 avdd.n128 avdd.n62 321.882
R10236 avdd.n114 avdd.n113 321.882
R10237 avdd.n60 avdd.n58 321.882
R10238 avdd.n76 avdd.n70 321.882
R10239 avdd.n93 avdd.n70 321.882
R10240 avdd.n93 avdd.n67 321.882
R10241 avdd.n97 avdd.n67 321.882
R10242 avdd.n98 avdd.n97 321.882
R10243 avdd.n98 avdd.n66 321.882
R10244 avdd.n102 avdd.n66 321.882
R10245 avdd.n646 avdd.n343 321.882
R10246 avdd.n632 avdd.n631 321.882
R10247 avdd.n341 avdd.n339 321.882
R10248 avdd.n618 avdd.n351 321.882
R10249 avdd.n604 avdd.n603 321.882
R10250 avdd.n349 avdd.n347 321.882
R10251 avdd.n590 avdd.n359 321.882
R10252 avdd.n576 avdd.n575 321.882
R10253 avdd.n357 avdd.n355 321.882
R10254 avdd.n562 avdd.n367 321.882
R10255 avdd.n548 avdd.n547 321.882
R10256 avdd.n365 avdd.n363 321.882
R10257 avdd.n534 avdd.n375 321.882
R10258 avdd.n520 avdd.n519 321.882
R10259 avdd.n373 avdd.n371 321.882
R10260 avdd.n506 avdd.n383 321.882
R10261 avdd.n492 avdd.n491 321.882
R10262 avdd.n381 avdd.n379 321.882
R10263 avdd.n478 avdd.n391 321.882
R10264 avdd.n464 avdd.n463 321.882
R10265 avdd.n389 avdd.n387 321.882
R10266 avdd.n450 avdd.n399 321.882
R10267 avdd.n436 avdd.n435 321.882
R10268 avdd.n397 avdd.n395 321.882
R10269 avdd.n422 avdd.n406 321.882
R10270 avdd.n412 avdd.n411 321.882
R10271 avdd.n424 avdd.n403 321.882
R10272 avdd.n666 avdd.n665 321.882
R10273 avdd.n794 avdd.n778 321.882
R10274 avdd.n799 avdd.n798 321.882
R10275 avdd.n798 avdd.n777 321.882
R10276 avdd.n810 avdd.n769 321.882
R10277 avdd.n806 avdd.n769 321.882
R10278 avdd.n819 avdd.n758 321.882
R10279 avdd.n771 avdd.n758 321.882
R10280 avdd.n824 avdd.n823 321.882
R10281 avdd.n823 avdd.n757 321.882
R10282 avdd.n835 avdd.n749 321.882
R10283 avdd.n831 avdd.n749 321.882
R10284 avdd.n844 avdd.n738 321.882
R10285 avdd.n751 avdd.n738 321.882
R10286 avdd.n849 avdd.n848 321.882
R10287 avdd.n848 avdd.n737 321.882
R10288 avdd.n860 avdd.n729 321.882
R10289 avdd.n856 avdd.n729 321.882
R10290 avdd.n869 avdd.n718 321.882
R10291 avdd.n731 avdd.n718 321.882
R10292 avdd.n874 avdd.n873 321.882
R10293 avdd.n873 avdd.n717 321.882
R10294 avdd.n885 avdd.n709 321.882
R10295 avdd.n881 avdd.n709 321.882
R10296 avdd.n894 avdd.n698 321.882
R10297 avdd.n711 avdd.n698 321.882
R10298 avdd.n899 avdd.n898 321.882
R10299 avdd.n898 avdd.n697 321.882
R10300 avdd.n910 avdd.n690 321.882
R10301 avdd.n906 avdd.n690 321.882
R10302 avdd.n685 avdd.n684 321.882
R10303 avdd.n686 avdd.n685 321.882
R10304 avdd.n786 avdd.n785 318.757
R10305 avdd.n1017 avdd.n946 300.048
R10306 avdd.n1151 avdd.n946 300.048
R10307 avdd.n976 avdd.t84 291.911
R10308 avdd.n1147 avdd.t80 291.911
R10309 avdd.n1148 avdd.t342 289.247
R10310 avdd.n1152 avdd.n945 281.601
R10311 avdd.t346 avdd.t426 272.962
R10312 avdd.n327 avdd.n326 271.068
R10313 avdd.n299 avdd.n298 271.068
R10314 avdd.n271 avdd.n270 271.068
R10315 avdd.n243 avdd.n242 271.068
R10316 avdd.n215 avdd.n214 271.068
R10317 avdd.n187 avdd.n186 271.068
R10318 avdd.n159 avdd.n158 271.068
R10319 avdd.n131 avdd.n130 271.068
R10320 avdd.n649 avdd.n648 271.068
R10321 avdd.n621 avdd.n620 271.068
R10322 avdd.n593 avdd.n592 271.068
R10323 avdd.n565 avdd.n564 271.068
R10324 avdd.n537 avdd.n536 271.068
R10325 avdd.n509 avdd.n508 271.068
R10326 avdd.n481 avdd.n480 271.068
R10327 avdd.n453 avdd.n452 271.068
R10328 avdd.n669 avdd.n668 271.068
R10329 avdd.n1299 avdd.n1218 257.882
R10330 avdd.n1285 avdd.n1219 257.882
R10331 avdd.n1229 avdd.t50 255.679
R10332 avdd.t137 avdd.n1229 255.679
R10333 avdd.n673 avdd.t333 252.983
R10334 avdd.n789 avdd.t420 252.983
R10335 avdd.n782 avdd.t438 252.983
R10336 avdd.n802 avdd.t279 252.983
R10337 avdd.n814 avdd.t37 252.983
R10338 avdd.n762 avdd.t69 252.983
R10339 avdd.n827 avdd.t239 252.983
R10340 avdd.n839 avdd.t217 252.983
R10341 avdd.n742 avdd.t300 252.983
R10342 avdd.n852 avdd.t198 252.983
R10343 avdd.n864 avdd.t265 252.983
R10344 avdd.n722 avdd.t39 252.983
R10345 avdd.n877 avdd.t432 252.983
R10346 avdd.n889 avdd.t271 252.983
R10347 avdd.n702 avdd.t430 252.983
R10348 avdd.n902 avdd.t267 252.983
R10349 avdd.n913 avdd.t186 252.983
R10350 avdd.n1143 avdd.t14 251.292
R10351 avdd.n1143 avdd.t21 251.292
R10352 avdd.t334 avdd.t426 241.649
R10353 avdd.n1352 avdd.n1351 241.459
R10354 avdd.n1348 avdd.n681 240.66
R10355 avdd.n1348 avdd.n1347 240.66
R10356 avdd.n1351 avdd.n678 240.66
R10357 avdd.t52 avdd.t56 233.565
R10358 avdd.t56 avdd.t60 233.565
R10359 avdd.t60 avdd.t66 233.565
R10360 avdd.t66 avdd.t58 233.565
R10361 avdd.t62 avdd.t64 233.565
R10362 avdd.t64 avdd.t54 233.565
R10363 avdd.t54 avdd.t244 233.565
R10364 avdd.t244 avdd.t246 233.565
R10365 avdd.n1158 avdd.t341 232.686
R10366 avdd.n970 avdd.t53 231.989
R10367 avdd.n985 avdd.t247 231.989
R10368 avdd.n1159 avdd.t345 231.974
R10369 avdd.n1158 avdd.t343 231.974
R10370 avdd.t159 avdd.n1068 227.345
R10371 avdd.n1122 avdd.t82 227.345
R10372 avdd.n423 avdd.t255 217.947
R10373 avdd.n1287 avdd.t346 216.344
R10374 avdd.n1291 avdd.t131 211.924
R10375 avdd.n960 avdd.n959 204.31
R10376 avdd.n1129 avdd.n1128 204.31
R10377 avdd.n1070 avdd.n1069 204.31
R10378 avdd.n978 avdd.n977 204.294
R10379 avdd.n980 avdd.n979 204.294
R10380 avdd.n982 avdd.n981 204.294
R10381 avdd.n984 avdd.n983 204.294
R10382 avdd.n1274 avdd.n1214 203.672
R10383 avdd.n1292 avdd.n1282 203.672
R10384 avdd.n325 avdd.t328 197.562
R10385 avdd.n297 avdd.t189 197.562
R10386 avdd.n269 avdd.t10 197.562
R10387 avdd.n241 avdd.t330 197.562
R10388 avdd.n213 avdd.t282 197.562
R10389 avdd.n185 avdd.t253 197.562
R10390 avdd.n157 avdd.t248 197.562
R10391 avdd.n129 avdd.t303 197.562
R10392 avdd.n647 avdd.t276 197.562
R10393 avdd.n619 avdd.t191 197.562
R10394 avdd.n591 avdd.t305 197.562
R10395 avdd.n563 avdd.t294 197.562
R10396 avdd.n535 avdd.t183 197.562
R10397 avdd.n507 avdd.t370 197.562
R10398 avdd.n479 avdd.t292 197.562
R10399 avdd.n451 avdd.t307 197.562
R10400 avdd.n1288 avdd.n1219 196.142
R10401 avdd.t340 avdd.n1148 195.042
R10402 avdd.n76 avdd.t296 193.774
R10403 avdd.n324 avdd.n323 185
R10404 avdd.n325 avdd.n324 185
R10405 avdd.n7 avdd.n6 185
R10406 avdd.n319 avdd.n309 185
R10407 avdd.n318 avdd.n310 185
R10408 avdd.n4 avdd.n1 185
R10409 avdd.n328 avdd.n2 185
R10410 avdd.n296 avdd.n295 185
R10411 avdd.n297 avdd.n296 185
R10412 avdd.n15 avdd.n14 185
R10413 avdd.n291 avdd.n281 185
R10414 avdd.n290 avdd.n282 185
R10415 avdd.n12 avdd.n9 185
R10416 avdd.n300 avdd.n10 185
R10417 avdd.n268 avdd.n267 185
R10418 avdd.n269 avdd.n268 185
R10419 avdd.n23 avdd.n22 185
R10420 avdd.n263 avdd.n253 185
R10421 avdd.n262 avdd.n254 185
R10422 avdd.n20 avdd.n17 185
R10423 avdd.n272 avdd.n18 185
R10424 avdd.n240 avdd.n239 185
R10425 avdd.n241 avdd.n240 185
R10426 avdd.n31 avdd.n30 185
R10427 avdd.n235 avdd.n225 185
R10428 avdd.n234 avdd.n226 185
R10429 avdd.n28 avdd.n25 185
R10430 avdd.n244 avdd.n26 185
R10431 avdd.n212 avdd.n211 185
R10432 avdd.n213 avdd.n212 185
R10433 avdd.n39 avdd.n38 185
R10434 avdd.n207 avdd.n197 185
R10435 avdd.n206 avdd.n198 185
R10436 avdd.n36 avdd.n33 185
R10437 avdd.n216 avdd.n34 185
R10438 avdd.n184 avdd.n183 185
R10439 avdd.n185 avdd.n184 185
R10440 avdd.n47 avdd.n46 185
R10441 avdd.n179 avdd.n169 185
R10442 avdd.n178 avdd.n170 185
R10443 avdd.n44 avdd.n41 185
R10444 avdd.n188 avdd.n42 185
R10445 avdd.n156 avdd.n155 185
R10446 avdd.n157 avdd.n156 185
R10447 avdd.n55 avdd.n54 185
R10448 avdd.n151 avdd.n141 185
R10449 avdd.n150 avdd.n142 185
R10450 avdd.n52 avdd.n49 185
R10451 avdd.n160 avdd.n50 185
R10452 avdd.n128 avdd.n127 185
R10453 avdd.n129 avdd.n128 185
R10454 avdd.n63 avdd.n62 185
R10455 avdd.n123 avdd.n113 185
R10456 avdd.n122 avdd.n114 185
R10457 avdd.n60 avdd.n57 185
R10458 avdd.n132 avdd.n58 185
R10459 avdd.n77 avdd.n76 185
R10460 avdd.n71 avdd.n70 185
R10461 avdd.n70 avdd.n69 185
R10462 avdd.n93 avdd.n92 185
R10463 avdd.n94 avdd.n93 185
R10464 avdd.n72 avdd.n67 185
R10465 avdd.n95 avdd.n67 185
R10466 avdd.n97 avdd.n68 185
R10467 avdd.n97 avdd.n96 185
R10468 avdd.n98 avdd.n65 185
R10469 avdd.n99 avdd.n98 185
R10470 avdd.n104 avdd.n66 185
R10471 avdd.n100 avdd.n66 185
R10472 avdd.n103 avdd.n102 185
R10473 avdd.n102 avdd.n101 185
R10474 avdd.n646 avdd.n645 185
R10475 avdd.n647 avdd.n646 185
R10476 avdd.n344 avdd.n343 185
R10477 avdd.n641 avdd.n631 185
R10478 avdd.n640 avdd.n632 185
R10479 avdd.n341 avdd.n338 185
R10480 avdd.n650 avdd.n339 185
R10481 avdd.n618 avdd.n617 185
R10482 avdd.n619 avdd.n618 185
R10483 avdd.n352 avdd.n351 185
R10484 avdd.n613 avdd.n603 185
R10485 avdd.n612 avdd.n604 185
R10486 avdd.n349 avdd.n346 185
R10487 avdd.n622 avdd.n347 185
R10488 avdd.n590 avdd.n589 185
R10489 avdd.n591 avdd.n590 185
R10490 avdd.n360 avdd.n359 185
R10491 avdd.n585 avdd.n575 185
R10492 avdd.n584 avdd.n576 185
R10493 avdd.n357 avdd.n354 185
R10494 avdd.n594 avdd.n355 185
R10495 avdd.n562 avdd.n561 185
R10496 avdd.n563 avdd.n562 185
R10497 avdd.n368 avdd.n367 185
R10498 avdd.n557 avdd.n547 185
R10499 avdd.n556 avdd.n548 185
R10500 avdd.n365 avdd.n362 185
R10501 avdd.n566 avdd.n363 185
R10502 avdd.n534 avdd.n533 185
R10503 avdd.n535 avdd.n534 185
R10504 avdd.n376 avdd.n375 185
R10505 avdd.n529 avdd.n519 185
R10506 avdd.n528 avdd.n520 185
R10507 avdd.n373 avdd.n370 185
R10508 avdd.n538 avdd.n371 185
R10509 avdd.n506 avdd.n505 185
R10510 avdd.n507 avdd.n506 185
R10511 avdd.n384 avdd.n383 185
R10512 avdd.n501 avdd.n491 185
R10513 avdd.n500 avdd.n492 185
R10514 avdd.n381 avdd.n378 185
R10515 avdd.n510 avdd.n379 185
R10516 avdd.n478 avdd.n477 185
R10517 avdd.n479 avdd.n478 185
R10518 avdd.n392 avdd.n391 185
R10519 avdd.n473 avdd.n463 185
R10520 avdd.n472 avdd.n464 185
R10521 avdd.n389 avdd.n386 185
R10522 avdd.n482 avdd.n387 185
R10523 avdd.n450 avdd.n449 185
R10524 avdd.n451 avdd.n450 185
R10525 avdd.n400 avdd.n399 185
R10526 avdd.n445 avdd.n435 185
R10527 avdd.n444 avdd.n436 185
R10528 avdd.n397 avdd.n394 185
R10529 avdd.n454 avdd.n395 185
R10530 avdd.n422 avdd.n421 185
R10531 avdd.n423 avdd.n422 185
R10532 avdd.n407 avdd.n406 185
R10533 avdd.n413 avdd.n412 185
R10534 avdd.n411 avdd.n402 185
R10535 avdd.n426 avdd.n403 185
R10536 avdd.n425 avdd.n424 185
R10537 avdd.n424 avdd.n423 185
R10538 avdd.n666 avdd.n664 185
R10539 avdd.n667 avdd.n666 185
R10540 avdd.n670 avdd.n665 185
R10541 avdd.n911 avdd.n910 185
R10542 avdd.n910 avdd.n909 185
R10543 avdd.n690 avdd.n689 185
R10544 avdd.n908 avdd.n690 185
R10545 avdd.n906 avdd.n905 185
R10546 avdd.n907 avdd.n906 185
R10547 avdd.n900 avdd.n899 185
R10548 avdd.n899 avdd.n693 185
R10549 avdd.n898 avdd.n696 185
R10550 avdd.n898 avdd.n897 185
R10551 avdd.n699 avdd.n697 185
R10552 avdd.n896 avdd.n697 185
R10553 avdd.n894 avdd.n893 185
R10554 avdd.n895 avdd.n894 185
R10555 avdd.n892 avdd.n698 185
R10556 avdd.n710 avdd.n698 185
R10557 avdd.n711 avdd.n705 185
R10558 avdd.n712 avdd.n711 185
R10559 avdd.n886 avdd.n885 185
R10560 avdd.n885 avdd.n884 185
R10561 avdd.n709 avdd.n708 185
R10562 avdd.n883 avdd.n709 185
R10563 avdd.n881 avdd.n880 185
R10564 avdd.n882 avdd.n881 185
R10565 avdd.n875 avdd.n874 185
R10566 avdd.n874 avdd.n713 185
R10567 avdd.n873 avdd.n716 185
R10568 avdd.n873 avdd.n872 185
R10569 avdd.n719 avdd.n717 185
R10570 avdd.n871 avdd.n717 185
R10571 avdd.n869 avdd.n868 185
R10572 avdd.n870 avdd.n869 185
R10573 avdd.n867 avdd.n718 185
R10574 avdd.n730 avdd.n718 185
R10575 avdd.n731 avdd.n725 185
R10576 avdd.n732 avdd.n731 185
R10577 avdd.n861 avdd.n860 185
R10578 avdd.n860 avdd.n859 185
R10579 avdd.n729 avdd.n728 185
R10580 avdd.n858 avdd.n729 185
R10581 avdd.n856 avdd.n855 185
R10582 avdd.n857 avdd.n856 185
R10583 avdd.n850 avdd.n849 185
R10584 avdd.n849 avdd.n733 185
R10585 avdd.n848 avdd.n736 185
R10586 avdd.n848 avdd.n847 185
R10587 avdd.n739 avdd.n737 185
R10588 avdd.n846 avdd.n737 185
R10589 avdd.n844 avdd.n843 185
R10590 avdd.n845 avdd.n844 185
R10591 avdd.n842 avdd.n738 185
R10592 avdd.n750 avdd.n738 185
R10593 avdd.n751 avdd.n745 185
R10594 avdd.n752 avdd.n751 185
R10595 avdd.n836 avdd.n835 185
R10596 avdd.n835 avdd.n834 185
R10597 avdd.n749 avdd.n748 185
R10598 avdd.n833 avdd.n749 185
R10599 avdd.n831 avdd.n830 185
R10600 avdd.n832 avdd.n831 185
R10601 avdd.n825 avdd.n824 185
R10602 avdd.n824 avdd.n753 185
R10603 avdd.n823 avdd.n756 185
R10604 avdd.n823 avdd.n822 185
R10605 avdd.n759 avdd.n757 185
R10606 avdd.n821 avdd.n757 185
R10607 avdd.n819 avdd.n818 185
R10608 avdd.n820 avdd.n819 185
R10609 avdd.n817 avdd.n758 185
R10610 avdd.n770 avdd.n758 185
R10611 avdd.n771 avdd.n765 185
R10612 avdd.n772 avdd.n771 185
R10613 avdd.n811 avdd.n810 185
R10614 avdd.n810 avdd.n809 185
R10615 avdd.n769 avdd.n768 185
R10616 avdd.n808 avdd.n769 185
R10617 avdd.n806 avdd.n805 185
R10618 avdd.n807 avdd.n806 185
R10619 avdd.n800 avdd.n799 185
R10620 avdd.n799 avdd.n773 185
R10621 avdd.n798 avdd.n776 185
R10622 avdd.n798 avdd.n797 185
R10623 avdd.n779 avdd.n777 185
R10624 avdd.n796 avdd.n777 185
R10625 avdd.n794 avdd.n793 185
R10626 avdd.n795 avdd.n794 185
R10627 avdd.n792 avdd.n778 185
R10628 avdd.n918 avdd.n684 185
R10629 avdd.n917 avdd.n685 185
R10630 avdd.n691 avdd.n685 185
R10631 avdd.n916 avdd.n686 185
R10632 avdd.n692 avdd.n686 185
R10633 avdd.n692 avdd.n691 175.386
R10634 avdd.n908 avdd.n907 175.386
R10635 avdd.n897 avdd.n896 175.386
R10636 avdd.n712 avdd.n710 175.386
R10637 avdd.n883 avdd.n882 175.386
R10638 avdd.n872 avdd.n871 175.386
R10639 avdd.n732 avdd.n730 175.386
R10640 avdd.n858 avdd.n857 175.386
R10641 avdd.n847 avdd.n846 175.386
R10642 avdd.n752 avdd.n750 175.386
R10643 avdd.n833 avdd.n832 175.386
R10644 avdd.n822 avdd.n821 175.386
R10645 avdd.n772 avdd.n770 175.386
R10646 avdd.n808 avdd.n807 175.386
R10647 avdd.n797 avdd.n796 175.386
R10648 avdd.n909 avdd.t266 169.905
R10649 avdd.t429 avdd.n693 169.905
R10650 avdd.n895 avdd.t270 169.905
R10651 avdd.n884 avdd.t431 169.905
R10652 avdd.t38 avdd.n713 169.905
R10653 avdd.n870 avdd.t264 169.905
R10654 avdd.n859 avdd.t197 169.905
R10655 avdd.t299 avdd.n733 169.905
R10656 avdd.n845 avdd.t216 169.905
R10657 avdd.n834 avdd.t238 169.905
R10658 avdd.t68 avdd.n753 169.905
R10659 avdd.n820 avdd.t36 169.905
R10660 avdd.n809 avdd.t278 169.905
R10661 avdd.t437 avdd.n773 169.905
R10662 avdd.n795 avdd.t419 169.905
R10663 avdd.t204 avdd.n1284 167.023
R10664 avdd.n1292 avdd.n1291 165.936
R10665 avdd.t336 avdd.n1287 156.744
R10666 avdd.n1294 avdd.n1293 155.859
R10667 avdd.n1298 avdd.n1297 155.859
R10668 avdd.t132 avdd.t204 153.764
R10669 avdd.t132 avdd.t336 153.764
R10670 avdd.n313 avdd.n312 153.571
R10671 avdd.n285 avdd.n284 153.571
R10672 avdd.n257 avdd.n256 153.571
R10673 avdd.n229 avdd.n228 153.571
R10674 avdd.n201 avdd.n200 153.571
R10675 avdd.n173 avdd.n172 153.571
R10676 avdd.n145 avdd.n144 153.571
R10677 avdd.n117 avdd.n116 153.571
R10678 avdd.n84 avdd.n83 153.571
R10679 avdd.n635 avdd.n634 153.571
R10680 avdd.n607 avdd.n606 153.571
R10681 avdd.n579 avdd.n578 153.571
R10682 avdd.n551 avdd.n550 153.571
R10683 avdd.n523 avdd.n522 153.571
R10684 avdd.n495 avdd.n494 153.571
R10685 avdd.n467 avdd.n466 153.571
R10686 avdd.n439 avdd.n438 153.571
R10687 avdd.n410 avdd.n409 153.571
R10688 avdd.t385 avdd.n1334 149.893
R10689 avdd.n1336 avdd.t405 149.893
R10690 avdd.t442 avdd.n1349 149.893
R10691 avdd.n1350 avdd.t263 149.893
R10692 avdd.n1204 avdd.n1163 148.329
R10693 avdd.n1337 avdd.n1331 125.742
R10694 avdd.n1329 avdd.n1312 125.742
R10695 avdd.n94 avdd.n69 120.317
R10696 avdd.n96 avdd.n95 120.317
R10697 avdd.n100 avdd.n99 120.317
R10698 avdd.n101 avdd.n100 120.317
R10699 avdd.n423 avdd.t240 117.838
R10700 avdd.n1266 avdd.t338 116.822
R10701 avdd.t58 avdd.n989 116.782
R10702 avdd.n989 avdd.t62 116.782
R10703 avdd.t240 avdd.t242 112.624
R10704 avdd.t399 avdd.t385 110.959
R10705 avdd.t415 avdd.t399 110.959
R10706 avdd.t395 avdd.t415 110.959
R10707 avdd.t411 avdd.t395 110.959
R10708 avdd.t407 avdd.t411 110.959
R10709 avdd.t389 avdd.t407 110.959
R10710 avdd.t403 avdd.t389 110.959
R10711 avdd.t401 avdd.t387 110.959
R10712 avdd.t397 avdd.t401 110.959
R10713 avdd.t413 avdd.t397 110.959
R10714 avdd.t393 avdd.t413 110.959
R10715 avdd.t409 avdd.t393 110.959
R10716 avdd.t391 avdd.t409 110.959
R10717 avdd.t405 avdd.t391 110.959
R10718 avdd.t441 avdd.t442 110.959
R10719 avdd.t127 avdd.t441 110.959
R10720 avdd.t434 avdd.t127 110.959
R10721 avdd.t433 avdd.t434 110.959
R10722 avdd.t90 avdd.t433 110.959
R10723 avdd.t43 avdd.t90 110.959
R10724 avdd.t42 avdd.t43 110.959
R10725 avdd.t140 avdd.t42 110.959
R10726 avdd.t212 avdd.t140 110.959
R10727 avdd.t211 avdd.t212 110.959
R10728 avdd.t112 avdd.t211 110.959
R10729 avdd.t311 avdd.t112 110.959
R10730 avdd.t312 avdd.t311 110.959
R10731 avdd.t163 avdd.t312 110.959
R10732 avdd.t323 avdd.t163 110.959
R10733 avdd.t322 avdd.t323 110.959
R10734 avdd.t103 avdd.t322 110.959
R10735 avdd.t310 avdd.t103 110.959
R10736 avdd.t309 avdd.t310 110.959
R10737 avdd.t178 avdd.t309 110.959
R10738 avdd.t349 avdd.t178 110.959
R10739 avdd.t348 avdd.t349 110.959
R10740 avdd.t167 avdd.t348 110.959
R10741 avdd.t356 avdd.t167 110.959
R10742 avdd.t357 avdd.t356 110.959
R10743 avdd.t157 avdd.t357 110.959
R10744 avdd.t436 avdd.t157 110.959
R10745 avdd.t435 avdd.t436 110.959
R10746 avdd.t165 avdd.t435 110.959
R10747 avdd.t320 avdd.t165 110.959
R10748 avdd.t321 avdd.t320 110.959
R10749 avdd.t125 avdd.t321 110.959
R10750 avdd.t439 avdd.t125 110.959
R10751 avdd.t440 avdd.t439 110.959
R10752 avdd.t176 avdd.t440 110.959
R10753 avdd.t40 avdd.t176 110.959
R10754 avdd.t41 avdd.t40 110.959
R10755 avdd.t180 avdd.t41 110.959
R10756 avdd.t375 avdd.t180 110.959
R10757 avdd.t376 avdd.t375 110.959
R10758 avdd.t152 avdd.t376 110.959
R10759 avdd.t302 avdd.t152 110.959
R10760 avdd.t301 avdd.t302 110.959
R10761 avdd.t92 avdd.t301 110.959
R10762 avdd.t262 avdd.t92 110.959
R10763 avdd.t263 avdd.t262 110.959
R10764 avdd.n325 avdd.t381 106.817
R10765 avdd.n297 avdd.t325 106.817
R10766 avdd.n269 avdd.t351 106.817
R10767 avdd.n241 avdd.t373 106.817
R10768 avdd.n213 avdd.t272 106.817
R10769 avdd.n185 avdd.t316 106.817
R10770 avdd.n157 avdd.t286 106.817
R10771 avdd.n129 avdd.t377 106.817
R10772 avdd.n647 avdd.t313 106.817
R10773 avdd.n619 avdd.t6 106.817
R10774 avdd.n591 avdd.t0 106.817
R10775 avdd.n563 avdd.t74 106.817
R10776 avdd.n535 avdd.t195 106.817
R10777 avdd.n507 avdd.t290 106.817
R10778 avdd.n479 avdd.t258 106.817
R10779 avdd.n451 avdd.t251 106.817
R10780 avdd.t354 avdd.n94 106.531
R10781 avdd.n1153 avdd.n944 105.788
R10782 avdd.t381 avdd.t206 102.091
R10783 avdd.t325 avdd.t181 102.091
R10784 avdd.t351 avdd.t214 102.091
R10785 avdd.t373 avdd.t284 102.091
R10786 avdd.t272 avdd.t274 102.091
R10787 avdd.t316 avdd.t318 102.091
R10788 avdd.t286 avdd.t187 102.091
R10789 avdd.t377 avdd.t379 102.091
R10790 avdd.t313 avdd.t268 102.091
R10791 avdd.t6 avdd.t8 102.091
R10792 avdd.t0 avdd.t2 102.091
R10793 avdd.t74 avdd.t70 102.091
R10794 avdd.t195 avdd.t193 102.091
R10795 avdd.t290 avdd.t280 102.091
R10796 avdd.t258 avdd.t208 102.091
R10797 avdd.t251 avdd.t72 102.091
R10798 avdd.t296 avdd.n69 101.564
R10799 avdd.n1151 avdd.n1150 99.0123
R10800 avdd.n1017 avdd.n1016 99.0123
R10801 avdd.n101 avdd.t260 97.7578
R10802 avdd.t199 avdd.n1222 96.5971
R10803 avdd.n956 avdd.n945 94.1181
R10804 avdd.n1063 avdd.n955 94.1181
R10805 avdd.n1135 avdd.n964 91.1064
R10806 avdd.t122 avdd.t199 88.8801
R10807 avdd.n1062 avdd.n968 87.7182
R10808 avdd.n6 avdd.n3 86.068
R10809 avdd.n310 avdd.n5 86.068
R10810 avdd.n326 avdd.n2 86.068
R10811 avdd.n309 avdd.n3 86.068
R10812 avdd.n5 avdd.n4 86.068
R10813 avdd.n14 avdd.n11 86.068
R10814 avdd.n282 avdd.n13 86.068
R10815 avdd.n298 avdd.n10 86.068
R10816 avdd.n281 avdd.n11 86.068
R10817 avdd.n13 avdd.n12 86.068
R10818 avdd.n22 avdd.n19 86.068
R10819 avdd.n254 avdd.n21 86.068
R10820 avdd.n270 avdd.n18 86.068
R10821 avdd.n253 avdd.n19 86.068
R10822 avdd.n21 avdd.n20 86.068
R10823 avdd.n30 avdd.n27 86.068
R10824 avdd.n226 avdd.n29 86.068
R10825 avdd.n242 avdd.n26 86.068
R10826 avdd.n225 avdd.n27 86.068
R10827 avdd.n29 avdd.n28 86.068
R10828 avdd.n38 avdd.n35 86.068
R10829 avdd.n198 avdd.n37 86.068
R10830 avdd.n214 avdd.n34 86.068
R10831 avdd.n197 avdd.n35 86.068
R10832 avdd.n37 avdd.n36 86.068
R10833 avdd.n46 avdd.n43 86.068
R10834 avdd.n170 avdd.n45 86.068
R10835 avdd.n186 avdd.n42 86.068
R10836 avdd.n169 avdd.n43 86.068
R10837 avdd.n45 avdd.n44 86.068
R10838 avdd.n54 avdd.n51 86.068
R10839 avdd.n142 avdd.n53 86.068
R10840 avdd.n158 avdd.n50 86.068
R10841 avdd.n141 avdd.n51 86.068
R10842 avdd.n53 avdd.n52 86.068
R10843 avdd.n62 avdd.n59 86.068
R10844 avdd.n114 avdd.n61 86.068
R10845 avdd.n130 avdd.n58 86.068
R10846 avdd.n113 avdd.n59 86.068
R10847 avdd.n61 avdd.n60 86.068
R10848 avdd.n343 avdd.n340 86.068
R10849 avdd.n632 avdd.n342 86.068
R10850 avdd.n648 avdd.n339 86.068
R10851 avdd.n631 avdd.n340 86.068
R10852 avdd.n342 avdd.n341 86.068
R10853 avdd.n351 avdd.n348 86.068
R10854 avdd.n604 avdd.n350 86.068
R10855 avdd.n620 avdd.n347 86.068
R10856 avdd.n603 avdd.n348 86.068
R10857 avdd.n350 avdd.n349 86.068
R10858 avdd.n359 avdd.n356 86.068
R10859 avdd.n576 avdd.n358 86.068
R10860 avdd.n592 avdd.n355 86.068
R10861 avdd.n575 avdd.n356 86.068
R10862 avdd.n358 avdd.n357 86.068
R10863 avdd.n367 avdd.n364 86.068
R10864 avdd.n548 avdd.n366 86.068
R10865 avdd.n564 avdd.n363 86.068
R10866 avdd.n547 avdd.n364 86.068
R10867 avdd.n366 avdd.n365 86.068
R10868 avdd.n375 avdd.n372 86.068
R10869 avdd.n520 avdd.n374 86.068
R10870 avdd.n536 avdd.n371 86.068
R10871 avdd.n519 avdd.n372 86.068
R10872 avdd.n374 avdd.n373 86.068
R10873 avdd.n383 avdd.n380 86.068
R10874 avdd.n492 avdd.n382 86.068
R10875 avdd.n508 avdd.n379 86.068
R10876 avdd.n491 avdd.n380 86.068
R10877 avdd.n382 avdd.n381 86.068
R10878 avdd.n391 avdd.n388 86.068
R10879 avdd.n464 avdd.n390 86.068
R10880 avdd.n480 avdd.n387 86.068
R10881 avdd.n463 avdd.n388 86.068
R10882 avdd.n390 avdd.n389 86.068
R10883 avdd.n399 avdd.n396 86.068
R10884 avdd.n436 avdd.n398 86.068
R10885 avdd.n452 avdd.n395 86.068
R10886 avdd.n435 avdd.n396 86.068
R10887 avdd.n398 avdd.n397 86.068
R10888 avdd.n406 avdd.n404 86.068
R10889 avdd.n411 avdd.n405 86.068
R10890 avdd.n412 avdd.n404 86.068
R10891 avdd.n405 avdd.n403 86.068
R10892 avdd.n668 avdd.n665 86.068
R10893 avdd.n785 avdd.t419 82.3568
R10894 avdd.n96 avdd.t360 72.6918
R10895 avdd.n1152 avdd.n1151 71.5299
R10896 avdd.n1018 avdd.n1017 71.5299
R10897 avdd.n785 avdd.n778 68.6629
R10898 avdd.n1013 avdd.t221 65.941
R10899 avdd.n1013 avdd.t35 65.941
R10900 avdd.n1011 avdd.t233 65.941
R10901 avdd.n1011 avdd.t26 65.941
R10902 avdd.n1009 avdd.t218 65.941
R10903 avdd.n1009 avdd.t29 65.941
R10904 avdd.n1007 avdd.t227 65.941
R10905 avdd.n1007 avdd.t22 65.941
R10906 avdd.n1005 avdd.t32 65.941
R10907 avdd.n1005 avdd.t228 65.941
R10908 avdd.n1003 avdd.t15 65.941
R10909 avdd.n1003 avdd.t234 65.941
R10910 avdd.n1001 avdd.t23 65.941
R10911 avdd.n1001 avdd.t219 65.941
R10912 avdd.n999 avdd.t33 65.941
R10913 avdd.n999 avdd.t229 65.941
R10914 avdd.n997 avdd.t16 65.941
R10915 avdd.n997 avdd.t236 65.941
R10916 avdd.n1088 avdd.t30 65.941
R10917 avdd.n1088 avdd.t134 65.941
R10918 avdd.n1090 avdd.t24 65.941
R10919 avdd.n1090 avdd.t87 65.941
R10920 avdd.n1092 avdd.t27 65.941
R10921 avdd.n1092 avdd.t114 65.941
R10922 avdd.n1094 avdd.t18 65.941
R10923 avdd.n1094 avdd.t171 65.941
R10924 avdd.n1096 avdd.t224 65.941
R10925 avdd.n1096 avdd.t96 65.941
R10926 avdd.n1098 avdd.t230 65.941
R10927 avdd.n1098 avdd.t119 65.941
R10928 avdd.n1100 avdd.t237 65.941
R10929 avdd.n1100 avdd.t147 65.941
R10930 avdd.n1102 avdd.t226 65.941
R10931 avdd.n1102 avdd.t107 65.941
R10932 avdd.n1104 avdd.t232 65.941
R10933 avdd.n1104 avdd.t129 65.941
R10934 avdd.t110 avdd.n1056 65.941
R10935 avdd.n1056 avdd.t223 65.941
R10936 avdd.n1053 avdd.t161 65.941
R10937 avdd.n1053 avdd.t235 65.941
R10938 avdd.n1050 avdd.t85 65.941
R10939 avdd.n1050 avdd.t220 65.941
R10940 avdd.t145 avdd.n1045 65.941
R10941 avdd.n1045 avdd.t231 65.941
R10942 avdd.t169 avdd.n1042 65.941
R10943 avdd.n1042 avdd.t34 65.941
R10944 avdd.n1039 avdd.t94 65.941
R10945 avdd.n1039 avdd.t19 65.941
R10946 avdd.n1036 avdd.t117 65.941
R10947 avdd.n1036 avdd.t25 65.941
R10948 avdd.t174 avdd.n1031 65.941
R10949 avdd.n1031 avdd.t13 65.941
R10950 avdd.n1028 avdd.t105 65.941
R10951 avdd.n1028 avdd.t20 65.941
R10952 avdd.n1228 avdd.t5 59.3422
R10953 avdd.n1335 avdd.t403 55.4795
R10954 avdd.t387 avdd.n1335 55.4795
R10955 avdd.n1327 avdd.t406 54.6604
R10956 avdd.n1310 avdd.t386 54.6604
R10957 avdd.n1276 avdd.t200 53.8832
R10958 avdd.n1270 avdd.t337 53.8832
R10959 avdd.n1269 avdd.t205 53.8832
R10960 avdd.n1210 avdd.n1209 50.4475
R10961 avdd.n1251 avdd.t136 49.5908
R10962 avdd.n1235 avdd.t136 49.5908
R10963 avdd.n325 avdd.n3 49.4675
R10964 avdd.n325 avdd.n5 49.4675
R10965 avdd.n326 avdd.n325 49.4675
R10966 avdd.n297 avdd.n11 49.4675
R10967 avdd.n297 avdd.n13 49.4675
R10968 avdd.n298 avdd.n297 49.4675
R10969 avdd.n269 avdd.n19 49.4675
R10970 avdd.n269 avdd.n21 49.4675
R10971 avdd.n270 avdd.n269 49.4675
R10972 avdd.n241 avdd.n27 49.4675
R10973 avdd.n241 avdd.n29 49.4675
R10974 avdd.n242 avdd.n241 49.4675
R10975 avdd.n213 avdd.n35 49.4675
R10976 avdd.n213 avdd.n37 49.4675
R10977 avdd.n214 avdd.n213 49.4675
R10978 avdd.n185 avdd.n43 49.4675
R10979 avdd.n185 avdd.n45 49.4675
R10980 avdd.n186 avdd.n185 49.4675
R10981 avdd.n157 avdd.n51 49.4675
R10982 avdd.n157 avdd.n53 49.4675
R10983 avdd.n158 avdd.n157 49.4675
R10984 avdd.n129 avdd.n59 49.4675
R10985 avdd.n129 avdd.n61 49.4675
R10986 avdd.n130 avdd.n129 49.4675
R10987 avdd.n647 avdd.n340 49.4675
R10988 avdd.n647 avdd.n342 49.4675
R10989 avdd.n648 avdd.n647 49.4675
R10990 avdd.n619 avdd.n348 49.4675
R10991 avdd.n619 avdd.n350 49.4675
R10992 avdd.n620 avdd.n619 49.4675
R10993 avdd.n591 avdd.n356 49.4675
R10994 avdd.n591 avdd.n358 49.4675
R10995 avdd.n592 avdd.n591 49.4675
R10996 avdd.n563 avdd.n364 49.4675
R10997 avdd.n563 avdd.n366 49.4675
R10998 avdd.n564 avdd.n563 49.4675
R10999 avdd.n535 avdd.n372 49.4675
R11000 avdd.n535 avdd.n374 49.4675
R11001 avdd.n536 avdd.n535 49.4675
R11002 avdd.n507 avdd.n380 49.4675
R11003 avdd.n507 avdd.n382 49.4675
R11004 avdd.n508 avdd.n507 49.4675
R11005 avdd.n479 avdd.n388 49.4675
R11006 avdd.n479 avdd.n390 49.4675
R11007 avdd.n480 avdd.n479 49.4675
R11008 avdd.n451 avdd.n396 49.4675
R11009 avdd.n451 avdd.n398 49.4675
R11010 avdd.n452 avdd.n451 49.4675
R11011 avdd.n423 avdd.n404 49.4675
R11012 avdd.n423 avdd.n405 49.4675
R11013 avdd.n668 avdd.n667 49.4675
R11014 avdd.n1326 avdd.n1325 49.1214
R11015 avdd.n1324 avdd.n1323 49.1214
R11016 avdd.n1322 avdd.n1321 49.1214
R11017 avdd.n1320 avdd.n1319 49.1214
R11018 avdd.n1318 avdd.n1317 49.1214
R11019 avdd.n1316 avdd.n1315 49.1214
R11020 avdd.n1314 avdd.n1313 49.1214
R11021 avdd.n1278 avdd.n1277 48.3442
R11022 avdd.n1280 avdd.n1279 48.3442
R11023 avdd.n1240 avdd.n1239 48.2034
R11024 avdd.n1242 avdd.n1241 48.2034
R11025 avdd.n1248 avdd.n1247 48.2034
R11026 avdd.n1255 avdd.n1254 48.2034
R11027 avdd.n1257 avdd.n1256 48.2034
R11028 avdd.n1259 avdd.n1258 48.2034
R11029 avdd.n1237 avdd.t101 48.0365
R11030 avdd.n1260 avdd.t123 48.0365
R11031 avdd.n99 avdd.t360 47.6258
R11032 avdd.t4 avdd.t428 47.3674
R11033 avdd.t428 avdd.t78 47.3674
R11034 avdd.t78 avdd.t425 47.3674
R11035 avdd.t150 avdd.t425 47.3674
R11036 avdd.t142 avdd.t203 47.3674
R11037 avdd.t201 avdd.t142 47.3674
R11038 avdd.t5 avdd.t201 47.3674
R11039 avdd.n1153 avdd.n1152 47.0593
R11040 avdd.n1065 avdd.n1063 44.8005
R11041 avdd.n1125 avdd.n945 44.8005
R11042 avdd.n1195 avdd.n1194 44.0934
R11043 avdd.n1085 avdd.n1084 43.2946
R11044 avdd.n1222 avdd.t421 42.8436
R11045 avdd.n1244 avdd.n1243 42.4975
R11046 avdd.n1246 avdd.n1236 42.4505
R11047 avdd.n1194 avdd.n1193 39.3333
R11048 avdd.n1016 avdd.n1015 37.0005
R11049 avdd.n1150 avdd.n1149 37.0005
R11050 avdd.n323 avdd.n7 36.1417
R11051 avdd.n319 avdd.n7 36.1417
R11052 avdd.n319 avdd.n318 36.1417
R11053 avdd.n318 avdd.n1 36.1417
R11054 avdd.n328 avdd.n1 36.1417
R11055 avdd.n328 avdd.n327 36.1417
R11056 avdd.n295 avdd.n15 36.1417
R11057 avdd.n291 avdd.n15 36.1417
R11058 avdd.n291 avdd.n290 36.1417
R11059 avdd.n290 avdd.n9 36.1417
R11060 avdd.n300 avdd.n9 36.1417
R11061 avdd.n300 avdd.n299 36.1417
R11062 avdd.n267 avdd.n23 36.1417
R11063 avdd.n263 avdd.n23 36.1417
R11064 avdd.n263 avdd.n262 36.1417
R11065 avdd.n262 avdd.n17 36.1417
R11066 avdd.n272 avdd.n17 36.1417
R11067 avdd.n272 avdd.n271 36.1417
R11068 avdd.n239 avdd.n31 36.1417
R11069 avdd.n235 avdd.n31 36.1417
R11070 avdd.n235 avdd.n234 36.1417
R11071 avdd.n234 avdd.n25 36.1417
R11072 avdd.n244 avdd.n25 36.1417
R11073 avdd.n244 avdd.n243 36.1417
R11074 avdd.n211 avdd.n39 36.1417
R11075 avdd.n207 avdd.n39 36.1417
R11076 avdd.n207 avdd.n206 36.1417
R11077 avdd.n206 avdd.n33 36.1417
R11078 avdd.n216 avdd.n33 36.1417
R11079 avdd.n216 avdd.n215 36.1417
R11080 avdd.n183 avdd.n47 36.1417
R11081 avdd.n179 avdd.n47 36.1417
R11082 avdd.n179 avdd.n178 36.1417
R11083 avdd.n178 avdd.n41 36.1417
R11084 avdd.n188 avdd.n41 36.1417
R11085 avdd.n188 avdd.n187 36.1417
R11086 avdd.n155 avdd.n55 36.1417
R11087 avdd.n151 avdd.n55 36.1417
R11088 avdd.n151 avdd.n150 36.1417
R11089 avdd.n150 avdd.n49 36.1417
R11090 avdd.n160 avdd.n49 36.1417
R11091 avdd.n160 avdd.n159 36.1417
R11092 avdd.n127 avdd.n63 36.1417
R11093 avdd.n123 avdd.n63 36.1417
R11094 avdd.n123 avdd.n122 36.1417
R11095 avdd.n122 avdd.n57 36.1417
R11096 avdd.n132 avdd.n57 36.1417
R11097 avdd.n132 avdd.n131 36.1417
R11098 avdd.n77 avdd.n71 36.1417
R11099 avdd.n92 avdd.n71 36.1417
R11100 avdd.n92 avdd.n72 36.1417
R11101 avdd.n72 avdd.n68 36.1417
R11102 avdd.n68 avdd.n65 36.1417
R11103 avdd.n104 avdd.n65 36.1417
R11104 avdd.n104 avdd.n103 36.1417
R11105 avdd.n645 avdd.n344 36.1417
R11106 avdd.n641 avdd.n344 36.1417
R11107 avdd.n641 avdd.n640 36.1417
R11108 avdd.n640 avdd.n338 36.1417
R11109 avdd.n650 avdd.n338 36.1417
R11110 avdd.n650 avdd.n649 36.1417
R11111 avdd.n617 avdd.n352 36.1417
R11112 avdd.n613 avdd.n352 36.1417
R11113 avdd.n613 avdd.n612 36.1417
R11114 avdd.n612 avdd.n346 36.1417
R11115 avdd.n622 avdd.n346 36.1417
R11116 avdd.n622 avdd.n621 36.1417
R11117 avdd.n589 avdd.n360 36.1417
R11118 avdd.n585 avdd.n360 36.1417
R11119 avdd.n585 avdd.n584 36.1417
R11120 avdd.n584 avdd.n354 36.1417
R11121 avdd.n594 avdd.n354 36.1417
R11122 avdd.n594 avdd.n593 36.1417
R11123 avdd.n561 avdd.n368 36.1417
R11124 avdd.n557 avdd.n368 36.1417
R11125 avdd.n557 avdd.n556 36.1417
R11126 avdd.n556 avdd.n362 36.1417
R11127 avdd.n566 avdd.n362 36.1417
R11128 avdd.n566 avdd.n565 36.1417
R11129 avdd.n533 avdd.n376 36.1417
R11130 avdd.n529 avdd.n376 36.1417
R11131 avdd.n529 avdd.n528 36.1417
R11132 avdd.n528 avdd.n370 36.1417
R11133 avdd.n538 avdd.n370 36.1417
R11134 avdd.n538 avdd.n537 36.1417
R11135 avdd.n505 avdd.n384 36.1417
R11136 avdd.n501 avdd.n384 36.1417
R11137 avdd.n501 avdd.n500 36.1417
R11138 avdd.n500 avdd.n378 36.1417
R11139 avdd.n510 avdd.n378 36.1417
R11140 avdd.n510 avdd.n509 36.1417
R11141 avdd.n477 avdd.n392 36.1417
R11142 avdd.n473 avdd.n392 36.1417
R11143 avdd.n473 avdd.n472 36.1417
R11144 avdd.n472 avdd.n386 36.1417
R11145 avdd.n482 avdd.n386 36.1417
R11146 avdd.n482 avdd.n481 36.1417
R11147 avdd.n449 avdd.n400 36.1417
R11148 avdd.n445 avdd.n400 36.1417
R11149 avdd.n445 avdd.n444 36.1417
R11150 avdd.n444 avdd.n394 36.1417
R11151 avdd.n454 avdd.n394 36.1417
R11152 avdd.n454 avdd.n453 36.1417
R11153 avdd.n421 avdd.n407 36.1417
R11154 avdd.n413 avdd.n407 36.1417
R11155 avdd.n413 avdd.n402 36.1417
R11156 avdd.n426 avdd.n402 36.1417
R11157 avdd.n426 avdd.n425 36.1417
R11158 avdd.n670 avdd.n664 36.1417
R11159 avdd.n670 avdd.n669 36.1417
R11160 avdd.n793 avdd.n792 36.1417
R11161 avdd.n792 avdd.n786 36.1417
R11162 avdd.n800 avdd.n776 36.1417
R11163 avdd.n779 avdd.n776 36.1417
R11164 avdd.n811 avdd.n768 36.1417
R11165 avdd.n805 avdd.n768 36.1417
R11166 avdd.n818 avdd.n817 36.1417
R11167 avdd.n817 avdd.n765 36.1417
R11168 avdd.n825 avdd.n756 36.1417
R11169 avdd.n759 avdd.n756 36.1417
R11170 avdd.n836 avdd.n748 36.1417
R11171 avdd.n830 avdd.n748 36.1417
R11172 avdd.n843 avdd.n842 36.1417
R11173 avdd.n842 avdd.n745 36.1417
R11174 avdd.n850 avdd.n736 36.1417
R11175 avdd.n739 avdd.n736 36.1417
R11176 avdd.n861 avdd.n728 36.1417
R11177 avdd.n855 avdd.n728 36.1417
R11178 avdd.n868 avdd.n867 36.1417
R11179 avdd.n867 avdd.n725 36.1417
R11180 avdd.n875 avdd.n716 36.1417
R11181 avdd.n719 avdd.n716 36.1417
R11182 avdd.n886 avdd.n708 36.1417
R11183 avdd.n880 avdd.n708 36.1417
R11184 avdd.n893 avdd.n892 36.1417
R11185 avdd.n892 avdd.n705 36.1417
R11186 avdd.n900 avdd.n696 36.1417
R11187 avdd.n699 avdd.n696 36.1417
R11188 avdd.n911 avdd.n689 36.1417
R11189 avdd.n905 avdd.n689 36.1417
R11190 avdd.n918 avdd.n917 36.1417
R11191 avdd.n917 avdd.n916 36.1417
R11192 avdd.t338 avdd.t122 32.9977
R11193 avdd.n1274 avdd.n1218 31.624
R11194 avdd.n1285 avdd.n1282 31.624
R11195 avdd.n1304 avdd.n1213 31.624
R11196 avdd.n987 avdd.n986 31.2476
R11197 avdd.n992 avdd.n991 31.2476
R11198 avdd.n955 avdd.n954 30.8338
R11199 avdd.n976 avdd.n954 30.8338
R11200 avdd.n956 avdd.n950 30.8338
R11201 avdd.n1147 avdd.n950 30.8338
R11202 avdd.n988 avdd.n987 30.8338
R11203 avdd.n991 avdd.n990 30.8338
R11204 avdd.n989 avdd.n976 28.7976
R11205 avdd.n1148 avdd.n1147 28.7976
R11206 avdd.n1195 avdd.n1190 28.3603
R11207 avdd.n1175 avdd.n1173 27.938
R11208 avdd.n959 avdd.t28 27.6955
R11209 avdd.n959 avdd.t225 27.6955
R11210 avdd.n1128 avdd.t222 27.6955
R11211 avdd.n1128 avdd.t81 27.6955
R11212 avdd.n1069 avdd.t159 27.6955
R11213 avdd.n1069 avdd.t31 27.6955
R11214 avdd.n977 avdd.t57 27.6955
R11215 avdd.n977 avdd.t61 27.6955
R11216 avdd.n979 avdd.t67 27.6955
R11217 avdd.n979 avdd.t59 27.6955
R11218 avdd.n981 avdd.t63 27.6955
R11219 avdd.n981 avdd.t65 27.6955
R11220 avdd.n983 avdd.t55 27.6955
R11221 avdd.n983 avdd.t245 27.6955
R11222 avdd.n1237 avdd.t98 25.5567
R11223 avdd.n1260 avdd.t121 25.5567
R11224 avdd.n1244 avdd.t153 25.4942
R11225 avdd.t203 avdd.t423 25.0145
R11226 avdd.n312 avdd.t383 23.5572
R11227 avdd.n284 avdd.t327 23.5572
R11228 avdd.n256 avdd.t353 23.5572
R11229 avdd.n228 avdd.t372 23.5572
R11230 avdd.n200 avdd.t275 23.5572
R11231 avdd.n172 avdd.t319 23.5572
R11232 avdd.n144 avdd.t288 23.5572
R11233 avdd.n116 avdd.t380 23.5572
R11234 avdd.n83 avdd.t361 23.5572
R11235 avdd.n634 avdd.t315 23.5572
R11236 avdd.n606 avdd.t9 23.5572
R11237 avdd.n578 avdd.t3 23.5572
R11238 avdd.n550 avdd.t76 23.5572
R11239 avdd.n522 avdd.t194 23.5572
R11240 avdd.n494 avdd.t289 23.5572
R11241 avdd.n466 avdd.t257 23.5572
R11242 avdd.n438 avdd.t250 23.5572
R11243 avdd.n409 avdd.t243 23.5572
R11244 avdd.t150 avdd.t423 22.3534
R11245 avdd.n74 avdd 20.0709
R11246 avdd.n1175 avdd.n1161 19.7066
R11247 avdd.n80 avdd 18.3657
R11248 avdd.n312 avdd.t207 17.8272
R11249 avdd.n284 avdd.t182 17.8272
R11250 avdd.n256 avdd.t215 17.8272
R11251 avdd.n228 avdd.t285 17.8272
R11252 avdd.n200 avdd.t350 17.8272
R11253 avdd.n172 avdd.t324 17.8272
R11254 avdd.n144 avdd.t188 17.8272
R11255 avdd.n116 avdd.t384 17.8272
R11256 avdd.n83 avdd.t355 17.8272
R11257 avdd.n634 avdd.t269 17.8272
R11258 avdd.n606 avdd.t418 17.8272
R11259 avdd.n578 avdd.t443 17.8272
R11260 avdd.n550 avdd.t71 17.8272
R11261 avdd.n522 avdd.t210 17.8272
R11262 avdd.n494 avdd.t281 17.8272
R11263 avdd.n466 avdd.t209 17.8272
R11264 avdd.n438 avdd.t73 17.8272
R11265 avdd.n409 avdd.t417 17.8272
R11266 avdd.n1205 avdd.n1162 17.7606
R11267 avdd.n336 avdd.n335 17.7258
R11268 avdd.n308 avdd.n307 17.7258
R11269 avdd.n280 avdd.n279 17.7258
R11270 avdd.n252 avdd.n251 17.7258
R11271 avdd.n224 avdd.n223 17.7258
R11272 avdd.n196 avdd.n195 17.7258
R11273 avdd.n168 avdd.n167 17.7258
R11274 avdd.n140 avdd.n139 17.7258
R11275 avdd.n112 avdd.n111 17.7258
R11276 avdd.n658 avdd.n657 17.7258
R11277 avdd.n630 avdd.n629 17.7258
R11278 avdd.n602 avdd.n601 17.7258
R11279 avdd.n574 avdd.n573 17.7258
R11280 avdd.n546 avdd.n545 17.7258
R11281 avdd.n518 avdd.n517 17.7258
R11282 avdd.n490 avdd.n489 17.7258
R11283 avdd.n462 avdd.n461 17.7258
R11284 avdd.n434 avdd.n433 17.7258
R11285 avdd.n1191 avdd.n1162 17.7066
R11286 avdd.n80 avdd.n79 17.3701
R11287 avdd.n79 avdd.n73 17.3701
R11288 avdd.t421 avdd.t4 16.4991
R11289 avdd.n1275 avdd.n1274 14.9605
R11290 avdd.n1282 avdd.n1281 14.9605
R11291 avdd.n1262 avdd.n1227 14.7677
R11292 avdd.n1189 avdd.n1170 14.6829
R11293 avdd.n1234 avdd.n1233 14.6449
R11294 avdd.n1068 avdd.t158 14.6083
R11295 avdd.n1122 avdd.t79 14.6083
R11296 avdd.n1262 avdd.n1253 14.5307
R11297 avdd.n1252 avdd.n1233 14.4078
R11298 avdd.n1187 avdd.n661 14.2404
R11299 avdd.n1289 avdd.n1288 14.2313
R11300 avdd.t132 avdd.n1289 14.2313
R11301 avdd.n1291 avdd.n1290 14.2313
R11302 avdd.n1290 avdd.t132 14.2313
R11303 avdd.n986 avdd.n985 14.0622
R11304 avdd.n1354 avdd.n1353 13.8347
R11305 avdd.n1344 avdd.n1343 13.8322
R11306 avdd.n936 avdd.n935 13.822
R11307 avdd.n1346 avdd.n937 13.822
R11308 avdd.n1066 avdd.n1065 13.8005
R11309 avdd.n1064 avdd.n966 13.8005
R11310 avdd.n996 avdd.n953 13.8005
R11311 avdd.n1127 avdd.n1126 13.8005
R11312 avdd.n1125 avdd.n1124 13.8005
R11313 avdd.n993 avdd.n992 13.8005
R11314 avdd.n95 avdd.t354 13.7868
R11315 avdd.n1188 avdd.n1172 13.5534
R11316 avdd.n1075 avdd.n1074 13.177
R11317 avdd.n1057 avdd.t109 12.679
R11318 avdd.n1052 avdd.t160 12.679
R11319 avdd.n1049 avdd.t83 12.679
R11320 avdd.n1046 avdd.t144 12.679
R11321 avdd.n1043 avdd.t168 12.679
R11322 avdd.n1038 avdd.t93 12.679
R11323 avdd.n1035 avdd.t116 12.679
R11324 avdd.n1032 avdd.t173 12.679
R11325 avdd.n1027 avdd.t104 12.679
R11326 avdd.n940 avdd.t133 12.679
R11327 avdd.n1106 avdd.t86 12.679
R11328 avdd.n1108 avdd.t113 12.679
R11329 avdd.n1110 avdd.t170 12.679
R11330 avdd.n1112 avdd.t95 12.679
R11331 avdd.n1114 avdd.t118 12.679
R11332 avdd.n1116 avdd.t146 12.679
R11333 avdd.n1118 avdd.t106 12.679
R11334 avdd.n1120 avdd.t128 12.679
R11335 avdd.n335 avdd.n334 12.541
R11336 avdd.n307 avdd.n306 12.541
R11337 avdd.n279 avdd.n278 12.541
R11338 avdd.n251 avdd.n250 12.541
R11339 avdd.n223 avdd.n222 12.541
R11340 avdd.n195 avdd.n194 12.541
R11341 avdd.n167 avdd.n166 12.541
R11342 avdd.n139 avdd.n138 12.541
R11343 avdd.n111 avdd.n110 12.541
R11344 avdd.n657 avdd.n656 12.541
R11345 avdd.n629 avdd.n628 12.541
R11346 avdd.n601 avdd.n600 12.541
R11347 avdd.n573 avdd.n572 12.541
R11348 avdd.n545 avdd.n544 12.541
R11349 avdd.n517 avdd.n516 12.541
R11350 avdd.n489 avdd.n488 12.541
R11351 avdd.n461 avdd.n460 12.541
R11352 avdd.n433 avdd.n432 12.541
R11353 avdd.n327 avdd 12.424
R11354 avdd.n299 avdd 12.424
R11355 avdd.n271 avdd 12.424
R11356 avdd.n243 avdd 12.424
R11357 avdd.n215 avdd 12.424
R11358 avdd.n187 avdd 12.424
R11359 avdd.n159 avdd 12.424
R11360 avdd.n131 avdd 12.424
R11361 avdd.n103 avdd 12.424
R11362 avdd.n649 avdd 12.424
R11363 avdd.n621 avdd 12.424
R11364 avdd.n593 avdd 12.424
R11365 avdd.n565 avdd 12.424
R11366 avdd.n537 avdd 12.424
R11367 avdd.n509 avdd 12.424
R11368 avdd.n481 avdd 12.424
R11369 avdd.n453 avdd 12.424
R11370 avdd.n425 avdd 12.424
R11371 avdd.n1186 avdd.n1173 12.2032
R11372 avdd.n1232 avdd.n1231 11.0005
R11373 avdd.n1264 avdd.n1263 11.0005
R11374 avdd.n1337 avdd.n1336 10.8829
R11375 avdd.n1334 avdd.n1329 10.8829
R11376 avdd.n1349 avdd.n1348 10.8829
R11377 avdd.n1351 avdd.n1350 10.8829
R11378 avdd.n1072 avdd.n1071 10.313
R11379 avdd.n1138 avdd.n961 10.313
R11380 avdd.n1132 avdd.n1131 10.313
R11381 avdd.n1284 avdd.n1283 10.2783
R11382 avdd.n1286 avdd.n1285 10.2783
R11383 avdd.n1287 avdd.n1286 10.2783
R11384 avdd.n1221 avdd.n1218 10.2783
R11385 avdd.n1222 avdd.n1221 10.2783
R11386 avdd.n1216 avdd.n1213 10.2783
R11387 avdd.n1228 avdd.n1216 10.2783
R11388 avdd.n1231 avdd.n1230 10.2783
R11389 avdd.n1265 avdd.n1264 10.2783
R11390 avdd.n1266 avdd.n1265 10.2783
R11391 avdd.t260 avdd.t358 10.0269
R11392 avdd.n1140 avdd.n957 9.71534
R11393 avdd.n332 avdd.n331 9.5406
R11394 avdd.n304 avdd.n303 9.5406
R11395 avdd.n276 avdd.n275 9.5406
R11396 avdd.n248 avdd.n247 9.5406
R11397 avdd.n220 avdd.n219 9.5406
R11398 avdd.n192 avdd.n191 9.5406
R11399 avdd.n164 avdd.n163 9.5406
R11400 avdd.n136 avdd.n135 9.5406
R11401 avdd.n108 avdd.n107 9.5406
R11402 avdd.n654 avdd.n653 9.5406
R11403 avdd.n626 avdd.n625 9.5406
R11404 avdd.n598 avdd.n597 9.5406
R11405 avdd.n570 avdd.n569 9.5406
R11406 avdd.n542 avdd.n541 9.5406
R11407 avdd.n514 avdd.n513 9.5406
R11408 avdd.n486 avdd.n485 9.5406
R11409 avdd.n458 avdd.n457 9.5406
R11410 avdd.n430 avdd.n429 9.5406
R11411 avdd.n1190 avdd.n661 9.42955
R11412 avdd.n81 avdd.n73 9.3005
R11413 avdd.n109 avdd.n108 9.3005
R11414 avdd.n108 avdd.n106 9.3005
R11415 avdd.n137 avdd.n136 9.3005
R11416 avdd.n136 avdd.n134 9.3005
R11417 avdd.n165 avdd.n164 9.3005
R11418 avdd.n164 avdd.n162 9.3005
R11419 avdd.n193 avdd.n192 9.3005
R11420 avdd.n192 avdd.n190 9.3005
R11421 avdd.n221 avdd.n220 9.3005
R11422 avdd.n220 avdd.n218 9.3005
R11423 avdd.n249 avdd.n248 9.3005
R11424 avdd.n248 avdd.n246 9.3005
R11425 avdd.n277 avdd.n276 9.3005
R11426 avdd.n276 avdd.n274 9.3005
R11427 avdd.n305 avdd.n304 9.3005
R11428 avdd.n304 avdd.n302 9.3005
R11429 avdd.n333 avdd.n332 9.3005
R11430 avdd.n332 avdd.n330 9.3005
R11431 avdd.n81 avdd.n80 9.3005
R11432 avdd.n88 avdd.n87 9.3005
R11433 avdd.n89 avdd.n88 9.3005
R11434 avdd.n120 avdd.n119 9.3005
R11435 avdd.n119 avdd.n118 9.3005
R11436 avdd.n148 avdd.n147 9.3005
R11437 avdd.n147 avdd.n146 9.3005
R11438 avdd.n176 avdd.n175 9.3005
R11439 avdd.n175 avdd.n174 9.3005
R11440 avdd.n204 avdd.n203 9.3005
R11441 avdd.n203 avdd.n202 9.3005
R11442 avdd.n232 avdd.n231 9.3005
R11443 avdd.n231 avdd.n230 9.3005
R11444 avdd.n260 avdd.n259 9.3005
R11445 avdd.n259 avdd.n258 9.3005
R11446 avdd.n288 avdd.n287 9.3005
R11447 avdd.n287 avdd.n286 9.3005
R11448 avdd.n316 avdd.n315 9.3005
R11449 avdd.n315 avdd.n314 9.3005
R11450 avdd.n78 avdd.n77 9.3005
R11451 avdd.n82 avdd.n71 9.3005
R11452 avdd.n92 avdd.n91 9.3005
R11453 avdd.n90 avdd.n72 9.3005
R11454 avdd.n85 avdd.n68 9.3005
R11455 avdd.n86 avdd.n65 9.3005
R11456 avdd.n105 avdd.n104 9.3005
R11457 avdd.n103 avdd.n64 9.3005
R11458 avdd.n127 avdd.n126 9.3005
R11459 avdd.n125 avdd.n63 9.3005
R11460 avdd.n124 avdd.n123 9.3005
R11461 avdd.n122 avdd.n121 9.3005
R11462 avdd.n115 avdd.n57 9.3005
R11463 avdd.n133 avdd.n132 9.3005
R11464 avdd.n131 avdd.n56 9.3005
R11465 avdd.n155 avdd.n154 9.3005
R11466 avdd.n153 avdd.n55 9.3005
R11467 avdd.n152 avdd.n151 9.3005
R11468 avdd.n150 avdd.n149 9.3005
R11469 avdd.n143 avdd.n49 9.3005
R11470 avdd.n161 avdd.n160 9.3005
R11471 avdd.n159 avdd.n48 9.3005
R11472 avdd.n183 avdd.n182 9.3005
R11473 avdd.n181 avdd.n47 9.3005
R11474 avdd.n180 avdd.n179 9.3005
R11475 avdd.n178 avdd.n177 9.3005
R11476 avdd.n171 avdd.n41 9.3005
R11477 avdd.n189 avdd.n188 9.3005
R11478 avdd.n187 avdd.n40 9.3005
R11479 avdd.n211 avdd.n210 9.3005
R11480 avdd.n209 avdd.n39 9.3005
R11481 avdd.n208 avdd.n207 9.3005
R11482 avdd.n206 avdd.n205 9.3005
R11483 avdd.n199 avdd.n33 9.3005
R11484 avdd.n217 avdd.n216 9.3005
R11485 avdd.n215 avdd.n32 9.3005
R11486 avdd.n239 avdd.n238 9.3005
R11487 avdd.n237 avdd.n31 9.3005
R11488 avdd.n236 avdd.n235 9.3005
R11489 avdd.n234 avdd.n233 9.3005
R11490 avdd.n227 avdd.n25 9.3005
R11491 avdd.n245 avdd.n244 9.3005
R11492 avdd.n243 avdd.n24 9.3005
R11493 avdd.n267 avdd.n266 9.3005
R11494 avdd.n265 avdd.n23 9.3005
R11495 avdd.n264 avdd.n263 9.3005
R11496 avdd.n262 avdd.n261 9.3005
R11497 avdd.n255 avdd.n17 9.3005
R11498 avdd.n273 avdd.n272 9.3005
R11499 avdd.n271 avdd.n16 9.3005
R11500 avdd.n295 avdd.n294 9.3005
R11501 avdd.n293 avdd.n15 9.3005
R11502 avdd.n292 avdd.n291 9.3005
R11503 avdd.n290 avdd.n289 9.3005
R11504 avdd.n283 avdd.n9 9.3005
R11505 avdd.n301 avdd.n300 9.3005
R11506 avdd.n299 avdd.n8 9.3005
R11507 avdd.n323 avdd.n322 9.3005
R11508 avdd.n321 avdd.n7 9.3005
R11509 avdd.n320 avdd.n319 9.3005
R11510 avdd.n318 avdd.n317 9.3005
R11511 avdd.n311 avdd.n1 9.3005
R11512 avdd.n329 avdd.n328 9.3005
R11513 avdd.n327 avdd.n0 9.3005
R11514 avdd.n431 avdd.n430 9.3005
R11515 avdd.n430 avdd.n428 9.3005
R11516 avdd.n459 avdd.n458 9.3005
R11517 avdd.n458 avdd.n456 9.3005
R11518 avdd.n487 avdd.n486 9.3005
R11519 avdd.n486 avdd.n484 9.3005
R11520 avdd.n515 avdd.n514 9.3005
R11521 avdd.n514 avdd.n512 9.3005
R11522 avdd.n543 avdd.n542 9.3005
R11523 avdd.n542 avdd.n540 9.3005
R11524 avdd.n571 avdd.n570 9.3005
R11525 avdd.n570 avdd.n568 9.3005
R11526 avdd.n599 avdd.n598 9.3005
R11527 avdd.n598 avdd.n596 9.3005
R11528 avdd.n627 avdd.n626 9.3005
R11529 avdd.n626 avdd.n624 9.3005
R11530 avdd.n655 avdd.n654 9.3005
R11531 avdd.n654 avdd.n652 9.3005
R11532 avdd.n417 avdd.n416 9.3005
R11533 avdd.n418 avdd.n417 9.3005
R11534 avdd.n442 avdd.n441 9.3005
R11535 avdd.n441 avdd.n440 9.3005
R11536 avdd.n470 avdd.n469 9.3005
R11537 avdd.n469 avdd.n468 9.3005
R11538 avdd.n498 avdd.n497 9.3005
R11539 avdd.n497 avdd.n496 9.3005
R11540 avdd.n526 avdd.n525 9.3005
R11541 avdd.n525 avdd.n524 9.3005
R11542 avdd.n554 avdd.n553 9.3005
R11543 avdd.n553 avdd.n552 9.3005
R11544 avdd.n582 avdd.n581 9.3005
R11545 avdd.n581 avdd.n580 9.3005
R11546 avdd.n610 avdd.n609 9.3005
R11547 avdd.n609 avdd.n608 9.3005
R11548 avdd.n638 avdd.n637 9.3005
R11549 avdd.n637 avdd.n636 9.3005
R11550 avdd.n421 avdd.n420 9.3005
R11551 avdd.n419 avdd.n407 9.3005
R11552 avdd.n414 avdd.n413 9.3005
R11553 avdd.n415 avdd.n402 9.3005
R11554 avdd.n427 avdd.n426 9.3005
R11555 avdd.n425 avdd.n401 9.3005
R11556 avdd.n449 avdd.n448 9.3005
R11557 avdd.n447 avdd.n400 9.3005
R11558 avdd.n446 avdd.n445 9.3005
R11559 avdd.n444 avdd.n443 9.3005
R11560 avdd.n437 avdd.n394 9.3005
R11561 avdd.n455 avdd.n454 9.3005
R11562 avdd.n453 avdd.n393 9.3005
R11563 avdd.n477 avdd.n476 9.3005
R11564 avdd.n475 avdd.n392 9.3005
R11565 avdd.n474 avdd.n473 9.3005
R11566 avdd.n472 avdd.n471 9.3005
R11567 avdd.n465 avdd.n386 9.3005
R11568 avdd.n483 avdd.n482 9.3005
R11569 avdd.n481 avdd.n385 9.3005
R11570 avdd.n505 avdd.n504 9.3005
R11571 avdd.n503 avdd.n384 9.3005
R11572 avdd.n502 avdd.n501 9.3005
R11573 avdd.n500 avdd.n499 9.3005
R11574 avdd.n493 avdd.n378 9.3005
R11575 avdd.n511 avdd.n510 9.3005
R11576 avdd.n509 avdd.n377 9.3005
R11577 avdd.n533 avdd.n532 9.3005
R11578 avdd.n531 avdd.n376 9.3005
R11579 avdd.n530 avdd.n529 9.3005
R11580 avdd.n528 avdd.n527 9.3005
R11581 avdd.n521 avdd.n370 9.3005
R11582 avdd.n539 avdd.n538 9.3005
R11583 avdd.n537 avdd.n369 9.3005
R11584 avdd.n561 avdd.n560 9.3005
R11585 avdd.n559 avdd.n368 9.3005
R11586 avdd.n558 avdd.n557 9.3005
R11587 avdd.n556 avdd.n555 9.3005
R11588 avdd.n549 avdd.n362 9.3005
R11589 avdd.n567 avdd.n566 9.3005
R11590 avdd.n565 avdd.n361 9.3005
R11591 avdd.n589 avdd.n588 9.3005
R11592 avdd.n587 avdd.n360 9.3005
R11593 avdd.n586 avdd.n585 9.3005
R11594 avdd.n584 avdd.n583 9.3005
R11595 avdd.n577 avdd.n354 9.3005
R11596 avdd.n595 avdd.n594 9.3005
R11597 avdd.n593 avdd.n353 9.3005
R11598 avdd.n617 avdd.n616 9.3005
R11599 avdd.n615 avdd.n352 9.3005
R11600 avdd.n614 avdd.n613 9.3005
R11601 avdd.n612 avdd.n611 9.3005
R11602 avdd.n605 avdd.n346 9.3005
R11603 avdd.n623 avdd.n622 9.3005
R11604 avdd.n621 avdd.n345 9.3005
R11605 avdd.n645 avdd.n644 9.3005
R11606 avdd.n643 avdd.n344 9.3005
R11607 avdd.n642 avdd.n641 9.3005
R11608 avdd.n640 avdd.n639 9.3005
R11609 avdd.n633 avdd.n338 9.3005
R11610 avdd.n651 avdd.n650 9.3005
R11611 avdd.n649 avdd.n337 9.3005
R11612 avdd.n1331 avdd.n1328 9.3005
R11613 avdd.n1340 avdd.n1312 9.3005
R11614 avdd.n673 avdd.n672 9.3005
R11615 avdd.n674 avdd.n673 9.3005
R11616 avdd.n664 avdd.n662 9.3005
R11617 avdd.n671 avdd.n670 9.3005
R11618 avdd.n669 avdd.n663 9.3005
R11619 avdd.n1305 avdd.n1304 9.3005
R11620 avdd.n1263 avdd.n1262 9.3005
R11621 avdd.n1233 avdd.n1232 9.3005
R11622 avdd.n1347 avdd.n1346 9.3005
R11623 avdd.n1344 avdd.n678 9.3005
R11624 avdd.n1353 avdd.n1352 9.3005
R11625 avdd.n935 avdd.n681 9.3005
R11626 avdd.n913 avdd.n687 9.3005
R11627 avdd.n914 avdd.n913 9.3005
R11628 avdd.n902 avdd.n694 9.3005
R11629 avdd.n903 avdd.n902 9.3005
R11630 avdd.n702 avdd.n701 9.3005
R11631 avdd.n703 avdd.n702 9.3005
R11632 avdd.n890 avdd.n889 9.3005
R11633 avdd.n889 avdd.n888 9.3005
R11634 avdd.n877 avdd.n714 9.3005
R11635 avdd.n878 avdd.n877 9.3005
R11636 avdd.n722 avdd.n721 9.3005
R11637 avdd.n723 avdd.n722 9.3005
R11638 avdd.n865 avdd.n864 9.3005
R11639 avdd.n864 avdd.n863 9.3005
R11640 avdd.n852 avdd.n734 9.3005
R11641 avdd.n853 avdd.n852 9.3005
R11642 avdd.n742 avdd.n741 9.3005
R11643 avdd.n743 avdd.n742 9.3005
R11644 avdd.n840 avdd.n839 9.3005
R11645 avdd.n839 avdd.n838 9.3005
R11646 avdd.n827 avdd.n754 9.3005
R11647 avdd.n828 avdd.n827 9.3005
R11648 avdd.n762 avdd.n761 9.3005
R11649 avdd.n763 avdd.n762 9.3005
R11650 avdd.n815 avdd.n814 9.3005
R11651 avdd.n814 avdd.n813 9.3005
R11652 avdd.n802 avdd.n774 9.3005
R11653 avdd.n803 avdd.n802 9.3005
R11654 avdd.n782 avdd.n781 9.3005
R11655 avdd.n783 avdd.n782 9.3005
R11656 avdd.n790 avdd.n789 9.3005
R11657 avdd.n789 avdd.n788 9.3005
R11658 avdd.n919 avdd.n918 9.3005
R11659 avdd.n917 avdd.n683 9.3005
R11660 avdd.n916 avdd.n915 9.3005
R11661 avdd.n912 avdd.n911 9.3005
R11662 avdd.n689 avdd.n688 9.3005
R11663 avdd.n905 avdd.n904 9.3005
R11664 avdd.n901 avdd.n900 9.3005
R11665 avdd.n696 avdd.n695 9.3005
R11666 avdd.n700 avdd.n699 9.3005
R11667 avdd.n893 avdd.n704 9.3005
R11668 avdd.n892 avdd.n891 9.3005
R11669 avdd.n706 avdd.n705 9.3005
R11670 avdd.n887 avdd.n886 9.3005
R11671 avdd.n708 avdd.n707 9.3005
R11672 avdd.n880 avdd.n879 9.3005
R11673 avdd.n876 avdd.n875 9.3005
R11674 avdd.n716 avdd.n715 9.3005
R11675 avdd.n720 avdd.n719 9.3005
R11676 avdd.n868 avdd.n724 9.3005
R11677 avdd.n867 avdd.n866 9.3005
R11678 avdd.n726 avdd.n725 9.3005
R11679 avdd.n862 avdd.n861 9.3005
R11680 avdd.n728 avdd.n727 9.3005
R11681 avdd.n855 avdd.n854 9.3005
R11682 avdd.n851 avdd.n850 9.3005
R11683 avdd.n736 avdd.n735 9.3005
R11684 avdd.n740 avdd.n739 9.3005
R11685 avdd.n843 avdd.n744 9.3005
R11686 avdd.n842 avdd.n841 9.3005
R11687 avdd.n746 avdd.n745 9.3005
R11688 avdd.n837 avdd.n836 9.3005
R11689 avdd.n748 avdd.n747 9.3005
R11690 avdd.n830 avdd.n829 9.3005
R11691 avdd.n826 avdd.n825 9.3005
R11692 avdd.n756 avdd.n755 9.3005
R11693 avdd.n760 avdd.n759 9.3005
R11694 avdd.n818 avdd.n764 9.3005
R11695 avdd.n817 avdd.n816 9.3005
R11696 avdd.n766 avdd.n765 9.3005
R11697 avdd.n812 avdd.n811 9.3005
R11698 avdd.n768 avdd.n767 9.3005
R11699 avdd.n805 avdd.n804 9.3005
R11700 avdd.n801 avdd.n800 9.3005
R11701 avdd.n776 avdd.n775 9.3005
R11702 avdd.n780 avdd.n779 9.3005
R11703 avdd.n793 avdd.n784 9.3005
R11704 avdd.n792 avdd.n791 9.3005
R11705 avdd.n787 avdd.n786 9.3005
R11706 avdd.n1345 avdd.n1344 9.2699
R11707 avdd.n1346 avdd.n1345 9.2699
R11708 avdd.n1207 avdd.n1206 8.56925
R11709 avdd.n948 avdd.n946 8.40959
R11710 avdd.n1148 avdd.n948 8.40959
R11711 avdd.n949 avdd.n947 8.40959
R11712 avdd.n1148 avdd.n949 8.40959
R11713 avdd.n1187 avdd.n1186 8.32145
R11714 avdd.n1309 avdd.n1308 7.90948
R11715 avdd.n1305 avdd.n1211 7.55653
R11716 avdd.n1268 avdd.n1211 7.55653
R11717 avdd.n1301 avdd.n1300 7.4005
R11718 avdd.t150 avdd.n1301 7.4005
R11719 avdd.n1303 avdd.n1302 7.4005
R11720 avdd.n1302 avdd.t150 7.4005
R11721 avdd.n1132 avdd.n1086 7.29542
R11722 avdd.n1309 avdd.n937 7.06613
R11723 avdd.n1268 avdd.n1212 7.06516
R11724 avdd.n1305 avdd.n1212 7.06516
R11725 avdd.n331 avdd 7.01471
R11726 avdd.n303 avdd 7.01471
R11727 avdd.n275 avdd 7.01471
R11728 avdd.n247 avdd 7.01471
R11729 avdd.n219 avdd 7.01471
R11730 avdd.n191 avdd 7.01471
R11731 avdd.n163 avdd 7.01471
R11732 avdd.n135 avdd 7.01471
R11733 avdd.n107 avdd 7.01471
R11734 avdd.n653 avdd 7.01471
R11735 avdd.n625 avdd 7.01471
R11736 avdd.n597 avdd 7.01471
R11737 avdd.n569 avdd 7.01471
R11738 avdd.n541 avdd 7.01471
R11739 avdd.n513 avdd 7.01471
R11740 avdd.n485 avdd 7.01471
R11741 avdd.n457 avdd 7.01471
R11742 avdd.n429 avdd 7.01471
R11743 avdd.n1072 avdd.n961 6.77003
R11744 avdd.n1137 avdd.n962 6.77003
R11745 avdd.n1073 avdd.n962 6.68605
R11746 avdd.n1133 avdd.n1132 6.6255
R11747 avdd.n1133 avdd.n963 6.60988
R11748 avdd.n974 avdd.n972 6.60764
R11749 avdd.n989 avdd.n974 6.60764
R11750 avdd.n973 avdd.n971 6.60764
R11751 avdd.n989 avdd.n973 6.60764
R11752 avdd.n1136 avdd.n963 6.59816
R11753 avdd.n1073 avdd.n1072 6.54933
R11754 avdd.n1140 avdd.n958 6.47706
R11755 avdd.n1020 avdd.n969 6.47706
R11756 avdd.n1020 avdd.n942 6.47706
R11757 avdd.n1342 avdd.n1341 5.7183
R11758 avdd.n1238 avdd.n1237 5.70732
R11759 avdd.n1261 avdd.n1260 5.70732
R11760 avdd.n1245 avdd.n1244 5.70732
R11761 avdd.n1238 avdd.n1233 5.70369
R11762 avdd.n1328 avdd.n1327 5.70305
R11763 avdd.n1262 avdd.n1261 5.70274
R11764 avdd.n1269 avdd.n1268 5.70242
R11765 avdd.n408 avdd 5.69343
R11766 avdd.n1341 avdd.n1340 5.6605
R11767 avdd.n1306 avdd.n1305 5.6605
R11768 avdd.n1250 avdd.n1249 5.6605
R11769 avdd.n975 avdd.n968 5.60656
R11770 avdd.n976 avdd.n975 5.60656
R11771 avdd.n1146 avdd.n944 5.60656
R11772 avdd.n1147 avdd.n1146 5.60656
R11773 avdd.n1325 avdd.t410 5.5395
R11774 avdd.n1325 avdd.t392 5.5395
R11775 avdd.n1323 avdd.t414 5.5395
R11776 avdd.n1323 avdd.t394 5.5395
R11777 avdd.n1321 avdd.t402 5.5395
R11778 avdd.n1321 avdd.t398 5.5395
R11779 avdd.n1319 avdd.t404 5.5395
R11780 avdd.n1319 avdd.t388 5.5395
R11781 avdd.n1317 avdd.t408 5.5395
R11782 avdd.n1317 avdd.t390 5.5395
R11783 avdd.n1315 avdd.t396 5.5395
R11784 avdd.n1315 avdd.t412 5.5395
R11785 avdd.n1313 avdd.t400 5.5395
R11786 avdd.n1313 avdd.t416 5.5395
R11787 avdd.n1246 avdd.t51 5.5395
R11788 avdd.t138 avdd.n1246 5.5395
R11789 avdd.n1209 avdd.t143 5.5395
R11790 avdd.n1209 avdd.t202 5.5395
R11791 avdd.n1277 avdd.t335 5.5395
R11792 avdd.n1277 avdd.t339 5.5395
R11793 avdd.n1279 avdd.t347 5.5395
R11794 avdd.n1279 avdd.t427 5.5395
R11795 avdd.n1243 avdd.t365 5.5395
R11796 avdd.n1243 avdd.t155 5.5395
R11797 avdd.n1239 avdd.t369 5.5395
R11798 avdd.n1239 avdd.t100 5.5395
R11799 avdd.t155 avdd.n1242 5.5395
R11800 avdd.n1242 avdd.t367 5.5395
R11801 avdd.n1247 avdd.t138 5.5395
R11802 avdd.n1247 avdd.t363 5.5395
R11803 avdd.n1254 avdd.t45 5.5395
R11804 avdd.n1254 avdd.t47 5.5395
R11805 avdd.n1256 avdd.t424 5.5395
R11806 avdd.n1256 avdd.t49 5.5395
R11807 avdd.t123 avdd.n1259 5.5395
R11808 avdd.n1259 avdd.t422 5.5395
R11809 avdd.n1339 avdd.n1328 5.48326
R11810 avdd.n1340 avdd.n1339 5.48326
R11811 avdd.n691 avdd.t185 5.48127
R11812 avdd.t266 avdd.n908 5.48127
R11813 avdd.n897 avdd.t429 5.48127
R11814 avdd.n710 avdd.t270 5.48127
R11815 avdd.t431 avdd.n883 5.48127
R11816 avdd.n872 avdd.t38 5.48127
R11817 avdd.n730 avdd.t264 5.48127
R11818 avdd.t197 avdd.n858 5.48127
R11819 avdd.n847 avdd.t299 5.48127
R11820 avdd.n750 avdd.t216 5.48127
R11821 avdd.t238 avdd.n833 5.48127
R11822 avdd.n822 avdd.t68 5.48127
R11823 avdd.n770 avdd.t36 5.48127
R11824 avdd.t278 avdd.n808 5.48127
R11825 avdd.n797 avdd.t437 5.48127
R11826 avdd.n1297 avdd.n1296 5.28621
R11827 avdd.n1296 avdd.t334 5.28621
R11828 avdd.n1295 avdd.n1294 5.28621
R11829 avdd.t334 avdd.n1295 5.28621
R11830 avdd.n1067 avdd.n957 5.22511
R11831 avdd.n1123 avdd.n943 5.22511
R11832 avdd.n1071 avdd.n1070 5.11573
R11833 avdd.t334 avdd.n1266 5.05652
R11834 avdd.n1178 avdd.n1177 4.89462
R11835 avdd.n1176 avdd.n1174 4.89462
R11836 avdd.n660 avdd.n659 4.7853
R11837 avdd.n1068 avdd.n1067 4.66083
R11838 avdd.n1123 avdd.n1122 4.66083
R11839 avdd.n1193 avdd.n1191 4.57145
R11840 avdd.n1160 avdd.n1159 4.54917
R11841 avdd.n1027 avdd.n967 4.5005
R11842 avdd.n1033 avdd.n1032 4.5005
R11843 avdd.n1035 avdd.n1034 4.5005
R11844 avdd.n1038 avdd.n1026 4.5005
R11845 avdd.n1044 avdd.n1043 4.5005
R11846 avdd.n1047 avdd.n1046 4.5005
R11847 avdd.n1049 avdd.n1048 4.5005
R11848 avdd.n1052 avdd.n995 4.5005
R11849 avdd.n1058 avdd.n1057 4.5005
R11850 avdd.n1138 avdd.n1137 4.5005
R11851 avdd.n1071 avdd.n962 4.5005
R11852 avdd.n1131 avdd.n963 4.5005
R11853 avdd.n1121 avdd.n1120 4.5005
R11854 avdd.n1119 avdd.n1118 4.5005
R11855 avdd.n1117 avdd.n1116 4.5005
R11856 avdd.n1115 avdd.n1114 4.5005
R11857 avdd.n1113 avdd.n1112 4.5005
R11858 avdd.n1111 avdd.n1110 4.5005
R11859 avdd.n1109 avdd.n1108 4.5005
R11860 avdd.n1107 avdd.n1106 4.5005
R11861 avdd.n941 avdd.n940 4.5005
R11862 avdd.n1130 avdd.n958 4.5005
R11863 avdd.n1140 avdd.n1139 4.5005
R11864 avdd.n1060 avdd.n1059 4.5005
R11865 avdd.n1024 avdd.n969 4.5005
R11866 avdd.n1021 avdd.n1020 4.5005
R11867 avdd.n1087 avdd.n942 4.5005
R11868 avdd.n1156 avdd.n1155 4.5005
R11869 avdd.n1308 avdd.n1207 4.4965
R11870 avdd.n80 avdd 4.46111
R11871 avdd.n80 avdd 4.46111
R11872 avdd.n1131 avdd.n1130 4.39112
R11873 avdd.n1076 avdd.n1075 4.30283
R11874 avdd.n1078 avdd.n1076 4.30283
R11875 avdd.n1077 avdd.n965 4.30283
R11876 avdd.n1081 avdd.n1077 4.30283
R11877 avdd.n994 avdd.n993 4.20743
R11878 avdd.n1338 avdd.n1330 4.20505
R11879 avdd.n1335 avdd.n1330 4.20505
R11880 avdd.n1333 avdd.n1332 4.20505
R11881 avdd.n1335 avdd.n1333 4.20505
R11882 avdd.n1139 avdd.n1138 4.16066
R11883 avdd.n1308 avdd.n1307 4.15861
R11884 avdd.n1307 avdd.n1306 4.01324
R11885 avdd.n1059 avdd.n994 3.98863
R11886 avdd.n1022 avdd.n1021 3.98863
R11887 avdd.n1087 avdd.n939 3.98863
R11888 avdd.n1024 avdd.n1023 3.98863
R11889 avdd.n1157 avdd.n1156 3.98863
R11890 avdd.n1340 avdd.n1311 3.91429
R11891 avdd.n1328 avdd.n1311 3.91429
R11892 avdd.n313 avdd 3.7406
R11893 avdd.n285 avdd 3.7406
R11894 avdd.n257 avdd 3.7406
R11895 avdd.n229 avdd 3.7406
R11896 avdd.n201 avdd 3.7406
R11897 avdd.n173 avdd 3.7406
R11898 avdd.n145 avdd 3.7406
R11899 avdd.n117 avdd 3.7406
R11900 avdd.n84 avdd 3.7406
R11901 avdd.n635 avdd 3.7406
R11902 avdd.n607 avdd 3.7406
R11903 avdd.n579 avdd 3.7406
R11904 avdd.n551 avdd 3.7406
R11905 avdd.n523 avdd 3.7406
R11906 avdd.n495 avdd 3.7406
R11907 avdd.n467 avdd 3.7406
R11908 avdd.n439 avdd 3.7406
R11909 avdd.n410 avdd 3.7406
R11910 avdd.n408 avdd 3.53935
R11911 avdd.n408 avdd 3.53935
R11912 avdd.n75 avdd 3.48691
R11913 avdd.n1185 avdd.n1184 3.24611
R11914 avdd.n1184 avdd.n1183 3.24611
R11915 avdd.n958 avdd.n943 3.23878
R11916 avdd.n1060 avdd.n969 3.23878
R11917 avdd.n1155 avdd.n942 3.23878
R11918 avdd.n1061 avdd.n957 3.14894
R11919 avdd.n1155 avdd.n1154 3.10206
R11920 avdd.n1154 avdd.n943 3.04738
R11921 avdd.n1061 avdd.n1060 3.01612
R11922 avdd.n659 avdd 2.67636
R11923 avdd.n1205 avdd.n1204 2.3255
R11924 avdd.n1206 avdd.n1205 2.307
R11925 avdd.n1180 avdd.n1172 2.17697
R11926 avdd.n1182 avdd.n1180 2.17697
R11927 avdd.n75 avdd 2.16773
R11928 avdd.n75 avdd 2.16773
R11929 avdd.n1307 avdd.n1208 1.97988
R11930 avdd.t48 avdd.n1228 1.86325
R11931 avdd.n1236 avdd.n1235 1.52433
R11932 avdd.n1134 avdd.n965 1.50638
R11933 avdd.n679 avdd.n677 1.4805
R11934 avdd.t167 avdd.n679 1.4805
R11935 avdd.n682 avdd.n680 1.4805
R11936 avdd.t167 avdd.n680 1.4805
R11937 avdd.n1251 avdd.n1250 1.31832
R11938 avdd.n935 avdd.n934 1.28283
R11939 avdd.n1019 avdd.n951 1.2505
R11940 avdd.n1143 avdd.n951 1.2505
R11941 avdd.n1144 avdd.n953 1.2505
R11942 avdd.n1144 avdd.n1143 1.2505
R11943 avdd.n1142 avdd.n1141 1.2505
R11944 avdd.n1143 avdd.n1142 1.2505
R11945 avdd.n1179 avdd.n1178 1.20965
R11946 avdd.n1181 avdd.n1179 1.20965
R11947 avdd.n936 avdd.n919 1.16964
R11948 avdd.n934 avdd.n933 1.15136
R11949 avdd.n933 avdd.n932 1.15136
R11950 avdd.n932 avdd.n931 1.15136
R11951 avdd.n931 avdd.n930 1.15136
R11952 avdd.n930 avdd.n929 1.15136
R11953 avdd.n929 avdd.n928 1.15136
R11954 avdd.n926 avdd.n925 1.15136
R11955 avdd.n925 avdd.n924 1.15136
R11956 avdd.n924 avdd.n923 1.15136
R11957 avdd.n923 avdd.n922 1.15136
R11958 avdd.n922 avdd.n921 1.15136
R11959 avdd.n921 avdd.n920 1.15136
R11960 avdd.n920 avdd.n676 1.15136
R11961 avdd.n1079 avdd.n964 1.14248
R11962 avdd.n1080 avdd.n1079 1.14248
R11963 avdd.n1084 avdd.n1083 1.14248
R11964 avdd.n1083 avdd.n1082 1.14248
R11965 avdd.n1197 avdd.n1196 1.14248
R11966 avdd.n1198 avdd.n1197 1.14248
R11967 avdd.n1353 avdd.n676 1.13628
R11968 avdd.n928 avdd.n927 1.0824
R11969 avdd.n1023 avdd.n1022 1.05355
R11970 avdd.n1022 avdd.n939 1.05355
R11971 avdd.n1225 avdd.n1223 1.03983
R11972 avdd.n1229 avdd.n1223 1.03983
R11973 avdd.n1226 avdd.n1224 1.03983
R11974 avdd.n1229 avdd.n1224 1.03983
R11975 avdd.n1164 avdd.n938 1.03383
R11976 avdd.n659 avdd 0.983
R11977 avdd.n1342 avdd.n1309 0.90425
R11978 avdd avdd.n661 0.876125
R11979 avdd.n1163 avdd.n1161 0.845955
R11980 avdd.n937 avdd.n936 0.83425
R11981 avdd.n1137 avdd.n1136 0.773938
R11982 avdd.n126 avdd 0.755
R11983 avdd.n154 avdd 0.755
R11984 avdd.n182 avdd 0.755
R11985 avdd.n210 avdd 0.755
R11986 avdd.n238 avdd 0.755
R11987 avdd.n266 avdd 0.755
R11988 avdd.n294 avdd 0.755
R11989 avdd.n322 avdd 0.755
R11990 avdd.n448 avdd 0.755
R11991 avdd.n476 avdd 0.755
R11992 avdd.n504 avdd 0.755
R11993 avdd.n532 avdd 0.755
R11994 avdd.n560 avdd 0.755
R11995 avdd.n588 avdd 0.755
R11996 avdd.n616 avdd 0.755
R11997 avdd.n644 avdd 0.755
R11998 avdd.n1130 avdd.n1129 0.725109
R11999 avdd.n1159 avdd.n1158 0.713391
R12000 avdd.n978 avdd.n970 0.695812
R12001 avdd.n980 avdd.n978 0.695812
R12002 avdd.n982 avdd.n980 0.695812
R12003 avdd.n984 avdd.n982 0.695812
R12004 avdd.n985 avdd.n984 0.695812
R12005 avdd.n1205 avdd.n1161 0.679554
R12006 avdd.n1139 avdd.n960 0.662609
R12007 avdd.n1355 avdd.n1354 0.624875
R12008 avdd.n78 avdd.n75 0.57
R12009 avdd.n660 avdd 0.563625
R12010 avdd.n1170 avdd.n1169 0.56281
R12011 avdd.n1169 avdd.n1168 0.56281
R12012 avdd.n1174 avdd.n1165 0.559412
R12013 avdd.n1167 avdd.n1165 0.559412
R12014 avdd.n1343 avdd.n675 0.55425
R12015 avdd.n1258 avdd.n1257 0.545446
R12016 avdd.n1257 avdd.n1255 0.545446
R12017 avdd.n1248 avdd.n1245 0.545446
R12018 avdd.n1241 avdd.n1240 0.545446
R12019 avdd.n1023 avdd.n994 0.527027
R12020 avdd.n1157 avdd.n939 0.527027
R12021 avdd.n75 avdd 0.51137
R12022 avdd.n1058 avdd.n995 0.486828
R12023 avdd.n1048 avdd.n995 0.486828
R12024 avdd.n1048 avdd.n1047 0.486828
R12025 avdd.n1047 avdd.n1044 0.486828
R12026 avdd.n1044 avdd.n1026 0.486828
R12027 avdd.n1034 avdd.n1026 0.486828
R12028 avdd.n1034 avdd.n1033 0.486828
R12029 avdd.n1033 avdd.n967 0.486828
R12030 avdd.n1014 avdd.n1012 0.486828
R12031 avdd.n1012 avdd.n1010 0.486828
R12032 avdd.n1010 avdd.n1008 0.486828
R12033 avdd.n1008 avdd.n1006 0.486828
R12034 avdd.n1006 avdd.n1004 0.486828
R12035 avdd.n1004 avdd.n1002 0.486828
R12036 avdd.n1002 avdd.n1000 0.486828
R12037 avdd.n1000 avdd.n998 0.486828
R12038 avdd.n1055 avdd.n1054 0.486828
R12039 avdd.n1054 avdd.n1051 0.486828
R12040 avdd.n1051 avdd.n1025 0.486828
R12041 avdd.n1041 avdd.n1025 0.486828
R12042 avdd.n1041 avdd.n1040 0.486828
R12043 avdd.n1040 avdd.n1037 0.486828
R12044 avdd.n1037 avdd.n1030 0.486828
R12045 avdd.n1030 avdd.n1029 0.486828
R12046 avdd.n1091 avdd.n1089 0.486828
R12047 avdd.n1093 avdd.n1091 0.486828
R12048 avdd.n1095 avdd.n1093 0.486828
R12049 avdd.n1097 avdd.n1095 0.486828
R12050 avdd.n1099 avdd.n1097 0.486828
R12051 avdd.n1101 avdd.n1099 0.486828
R12052 avdd.n1103 avdd.n1101 0.486828
R12053 avdd.n1105 avdd.n1103 0.486828
R12054 avdd.n1107 avdd.n941 0.486828
R12055 avdd.n1109 avdd.n1107 0.486828
R12056 avdd.n1111 avdd.n1109 0.486828
R12057 avdd.n1113 avdd.n1111 0.486828
R12058 avdd.n1115 avdd.n1113 0.486828
R12059 avdd.n1117 avdd.n1115 0.486828
R12060 avdd.n1119 avdd.n1117 0.486828
R12061 avdd.n1121 avdd.n1119 0.486828
R12062 avdd.n1066 avdd.n967 0.477062
R12063 avdd.n998 avdd.n996 0.477062
R12064 avdd.n1029 avdd.n966 0.477062
R12065 avdd.n1127 avdd.n1105 0.477062
R12066 avdd.n1124 avdd.n1121 0.477062
R12067 avdd.n1202 avdd.n1201 0.458421
R12068 avdd.n1201 avdd.n1200 0.458421
R12069 avdd.n1207 avdd.n938 0.4145
R12070 avdd.n661 avdd.n660 0.407375
R12071 avdd.n1059 avdd.n1058 0.340344
R12072 avdd.n1021 avdd.n1014 0.340344
R12073 avdd.n1055 avdd.n1024 0.340344
R12074 avdd.n1089 avdd.n1087 0.340344
R12075 avdd.n1156 avdd.n941 0.340344
R12076 avdd.n1355 avdd 0.32398
R12077 avdd.n1067 avdd.n1066 0.318859
R12078 avdd.n996 avdd.n960 0.318859
R12079 avdd.n1070 avdd.n966 0.318859
R12080 avdd.n1129 avdd.n1127 0.318859
R12081 avdd.n1124 avdd.n1123 0.318859
R12082 avdd.n1249 avdd.n1208 0.316162
R12083 avdd.n1171 avdd.n1166 0.306791
R12084 avdd.n1199 avdd.n1166 0.306791
R12085 avdd.n1280 avdd.n1278 0.291392
R12086 avdd.n1278 avdd.n1276 0.291392
R12087 avdd.n1235 avdd.n1234 0.284354
R12088 avdd.n1252 avdd.n1251 0.284354
R12089 avdd.n1354 avdd.n675 0.2805
R12090 avdd.n1249 avdd.n1248 0.273291
R12091 avdd.n1261 avdd.n1258 0.272973
R12092 avdd.n1245 avdd.n1241 0.272973
R12093 avdd.n1240 avdd.n1238 0.272973
R12094 avdd.n993 avdd.n970 0.262219
R12095 avdd avdd.n912 0.248811
R12096 avdd avdd.n901 0.248811
R12097 avdd.n704 avdd 0.248811
R12098 avdd avdd.n887 0.248811
R12099 avdd avdd.n876 0.248811
R12100 avdd.n724 avdd 0.248811
R12101 avdd avdd.n862 0.248811
R12102 avdd avdd.n851 0.248811
R12103 avdd.n744 avdd 0.248811
R12104 avdd avdd.n837 0.248811
R12105 avdd avdd.n826 0.248811
R12106 avdd.n764 avdd 0.248811
R12107 avdd avdd.n812 0.248811
R12108 avdd avdd.n801 0.248811
R12109 avdd.n784 avdd 0.248811
R12110 avdd.n1270 avdd.n1269 0.246297
R12111 avdd.n1134 avdd.n1133 0.245237
R12112 avdd.n1074 avdd.n1073 0.245237
R12113 avdd.n1206 avdd 0.242804
R12114 avdd.n1062 avdd.n1061 0.238962
R12115 avdd.n1154 avdd.n1153 0.238962
R12116 avdd.n1343 avdd.n1342 0.238625
R12117 avdd.n1255 avdd.n1208 0.229784
R12118 avdd.n1160 avdd.n1157 0.227878
R12119 avdd.n1332 avdd.n1311 0.227329
R12120 avdd.n1339 avdd.n1338 0.227329
R12121 avdd.n1281 avdd.n1280 0.1885
R12122 avdd.n1275 avdd.n1273 0.183736
R12123 avdd.n74 avdd 0.177503
R12124 avdd.n675 avdd.n674 0.175331
R12125 avdd.n1186 avdd.n1185 0.166571
R12126 avdd.n1306 avdd.n1210 0.156108
R12127 avdd.n1293 avdd.n1212 0.126176
R12128 avdd.n1298 avdd.n1211 0.126176
R12129 avdd.n1193 avdd.n1192 0.1245
R12130 avdd.n1234 avdd.n1227 0.123345
R12131 avdd.n1253 avdd.n1252 0.123345
R12132 avdd.n1188 avdd.n1187 0.113915
R12133 avdd.n1314 avdd.n1310 0.113554
R12134 avdd.n1316 avdd.n1314 0.113554
R12135 avdd.n1318 avdd.n1316 0.113554
R12136 avdd.n1320 avdd.n1318 0.113554
R12137 avdd.n1322 avdd.n1320 0.113554
R12138 avdd.n1324 avdd.n1322 0.113554
R12139 avdd.n1326 avdd.n1324 0.113554
R12140 avdd.n1327 avdd.n1326 0.113554
R12141 avdd.n1273 avdd.n1272 0.113554
R12142 avdd.n1272 avdd.n1271 0.113554
R12143 avdd.n1250 avdd.n1236 0.0934054
R12144 avdd avdd.n74 0.0845052
R12145 avdd.n671 avdd.n663 0.0815811
R12146 avdd.n919 avdd.n683 0.0815811
R12147 avdd.n912 avdd.n688 0.0815811
R12148 avdd.n901 avdd.n695 0.0815811
R12149 avdd.n891 avdd.n704 0.0815811
R12150 avdd.n887 avdd.n707 0.0815811
R12151 avdd.n876 avdd.n715 0.0815811
R12152 avdd.n866 avdd.n724 0.0815811
R12153 avdd.n862 avdd.n727 0.0815811
R12154 avdd.n851 avdd.n735 0.0815811
R12155 avdd.n841 avdd.n744 0.0815811
R12156 avdd.n837 avdd.n747 0.0815811
R12157 avdd.n826 avdd.n755 0.0815811
R12158 avdd.n816 avdd.n764 0.0815811
R12159 avdd.n812 avdd.n767 0.0815811
R12160 avdd.n801 avdd.n775 0.0815811
R12161 avdd.n791 avdd.n784 0.0815811
R12162 avdd.n1345 avdd.n682 0.0793136
R12163 avdd.n927 avdd.n677 0.0793136
R12164 avdd.n1086 avdd.n961 0.0766719
R12165 avdd.n927 avdd.n926 0.0694655
R12166 avdd.n1141 avdd.n1140 0.0674065
R12167 avdd.n1020 avdd.n1019 0.0674065
R12168 avdd.n1086 avdd.n1085 0.0650833
R12169 avdd.n1136 avdd.n1135 0.0650833
R12170 avdd.n1177 avdd.n1173 0.0641986
R12171 avdd.n1196 avdd.n1195 0.0608896
R12172 avdd.n315 avdd.n313 0.0579519
R12173 avdd.n287 avdd.n285 0.0579519
R12174 avdd.n259 avdd.n257 0.0579519
R12175 avdd.n231 avdd.n229 0.0579519
R12176 avdd.n203 avdd.n201 0.0579519
R12177 avdd.n175 avdd.n173 0.0579519
R12178 avdd.n147 avdd.n145 0.0579519
R12179 avdd.n119 avdd.n117 0.0579519
R12180 avdd.n88 avdd.n84 0.0579519
R12181 avdd.n637 avdd.n635 0.0579519
R12182 avdd.n609 avdd.n607 0.0579519
R12183 avdd.n581 avdd.n579 0.0579519
R12184 avdd.n553 avdd.n551 0.0579519
R12185 avdd.n525 avdd.n523 0.0579519
R12186 avdd.n497 avdd.n495 0.0579519
R12187 avdd.n469 avdd.n467 0.0579519
R12188 avdd.n441 avdd.n439 0.0579519
R12189 avdd.n417 avdd.n410 0.0579519
R12190 avdd.n1227 avdd.n1225 0.0558571
R12191 avdd.n1253 avdd.n1226 0.0558571
R12192 avdd.n672 avdd.n662 0.0553986
R12193 avdd.n915 avdd.n687 0.0553986
R12194 avdd.n904 avdd.n694 0.0553986
R12195 avdd.n701 avdd.n700 0.0553986
R12196 avdd.n890 avdd.n706 0.0553986
R12197 avdd.n879 avdd.n714 0.0553986
R12198 avdd.n721 avdd.n720 0.0553986
R12199 avdd.n865 avdd.n726 0.0553986
R12200 avdd.n854 avdd.n734 0.0553986
R12201 avdd.n741 avdd.n740 0.0553986
R12202 avdd.n840 avdd.n746 0.0553986
R12203 avdd.n829 avdd.n754 0.0553986
R12204 avdd.n761 avdd.n760 0.0553986
R12205 avdd.n815 avdd.n766 0.0553986
R12206 avdd.n804 avdd.n774 0.0553986
R12207 avdd.n781 avdd.n780 0.0553986
R12208 avdd.n790 avdd.n787 0.0553986
R12209 avdd avdd.n1355 0.04675
R12210 avdd.n1276 avdd.n1275 0.0436892
R12211 avdd.n1341 avdd.n1310 0.0430541
R12212 avdd.n1281 avdd.n1270 0.0430541
R12213 avdd.n663 avdd 0.0410405
R12214 avdd avdd.n90 0.04
R12215 avdd avdd.n124 0.04
R12216 avdd avdd.n152 0.04
R12217 avdd avdd.n180 0.04
R12218 avdd avdd.n208 0.04
R12219 avdd avdd.n236 0.04
R12220 avdd avdd.n264 0.04
R12221 avdd avdd.n292 0.04
R12222 avdd avdd.n320 0.04
R12223 avdd avdd.n419 0.04
R12224 avdd avdd.n446 0.04
R12225 avdd avdd.n474 0.04
R12226 avdd avdd.n502 0.04
R12227 avdd avdd.n530 0.04
R12228 avdd avdd.n558 0.04
R12229 avdd avdd.n586 0.04
R12230 avdd avdd.n614 0.04
R12231 avdd avdd.n642 0.04
R12232 avdd.n1191 avdd.n938 0.0375
R12233 avdd avdd.n86 0.0365
R12234 avdd avdd.n115 0.0365
R12235 avdd avdd.n143 0.0365
R12236 avdd avdd.n171 0.0365
R12237 avdd avdd.n199 0.0365
R12238 avdd avdd.n227 0.0365
R12239 avdd avdd.n255 0.0365
R12240 avdd avdd.n283 0.0365
R12241 avdd avdd.n311 0.0365
R12242 avdd avdd.n415 0.0365
R12243 avdd avdd.n437 0.0365
R12244 avdd avdd.n465 0.0365
R12245 avdd avdd.n493 0.0365
R12246 avdd avdd.n521 0.0365
R12247 avdd avdd.n549 0.0365
R12248 avdd avdd.n577 0.0365
R12249 avdd avdd.n605 0.0365
R12250 avdd avdd.n633 0.0365
R12251 avdd.n914 avdd 0.0351284
R12252 avdd.n903 avdd 0.0351284
R12253 avdd avdd.n703 0.0351284
R12254 avdd.n888 avdd 0.0351284
R12255 avdd.n878 avdd 0.0351284
R12256 avdd avdd.n723 0.0351284
R12257 avdd.n863 avdd 0.0351284
R12258 avdd.n853 avdd 0.0351284
R12259 avdd avdd.n743 0.0351284
R12260 avdd.n838 avdd 0.0351284
R12261 avdd.n828 avdd 0.0351284
R12262 avdd avdd.n763 0.0351284
R12263 avdd.n813 avdd 0.0351284
R12264 avdd.n803 avdd 0.0351284
R12265 avdd avdd.n783 0.0351284
R12266 avdd.n788 avdd 0.0351284
R12267 avdd.n1203 avdd.n1162 0.0324588
R12268 avdd.n106 avdd 0.032
R12269 avdd.n134 avdd 0.032
R12270 avdd.n162 avdd 0.032
R12271 avdd.n190 avdd 0.032
R12272 avdd.n218 avdd 0.032
R12273 avdd.n246 avdd 0.032
R12274 avdd.n274 avdd 0.032
R12275 avdd.n302 avdd 0.032
R12276 avdd.n330 avdd 0.032
R12277 avdd.n428 avdd 0.032
R12278 avdd.n456 avdd 0.032
R12279 avdd.n484 avdd 0.032
R12280 avdd.n512 avdd 0.032
R12281 avdd.n540 avdd 0.032
R12282 avdd.n568 avdd 0.032
R12283 avdd.n596 avdd 0.032
R12284 avdd.n624 avdd 0.032
R12285 avdd.n652 avdd 0.032
R12286 avdd.n1190 avdd.n1189 0.0301178
R12287 avdd.n1176 avdd.n1175 0.0300238
R12288 avdd.n1271 avdd.n1210 0.0287635
R12289 avdd.n81 avdd 0.028
R12290 avdd.n672 avdd.n671 0.0266824
R12291 avdd.n687 avdd.n683 0.0266824
R12292 avdd.n694 avdd.n688 0.0266824
R12293 avdd.n701 avdd.n695 0.0266824
R12294 avdd.n891 avdd.n890 0.0266824
R12295 avdd.n714 avdd.n707 0.0266824
R12296 avdd.n721 avdd.n715 0.0266824
R12297 avdd.n866 avdd.n865 0.0266824
R12298 avdd.n734 avdd.n727 0.0266824
R12299 avdd.n741 avdd.n735 0.0266824
R12300 avdd.n841 avdd.n840 0.0266824
R12301 avdd.n754 avdd.n747 0.0266824
R12302 avdd.n761 avdd.n755 0.0266824
R12303 avdd.n816 avdd.n815 0.0266824
R12304 avdd.n774 avdd.n767 0.0266824
R12305 avdd.n781 avdd.n775 0.0266824
R12306 avdd.n791 avdd.n790 0.0266824
R12307 avdd.n91 avdd 0.0245
R12308 avdd.n85 avdd 0.0245
R12309 avdd avdd.n125 0.0245
R12310 avdd.n121 avdd 0.0245
R12311 avdd avdd.n153 0.0245
R12312 avdd.n149 avdd 0.0245
R12313 avdd avdd.n181 0.0245
R12314 avdd.n177 avdd 0.0245
R12315 avdd avdd.n209 0.0245
R12316 avdd.n205 avdd 0.0245
R12317 avdd avdd.n237 0.0245
R12318 avdd.n233 avdd 0.0245
R12319 avdd avdd.n265 0.0245
R12320 avdd.n261 avdd 0.0245
R12321 avdd avdd.n293 0.0245
R12322 avdd.n289 avdd 0.0245
R12323 avdd avdd.n321 0.0245
R12324 avdd.n317 avdd 0.0245
R12325 avdd.n414 avdd 0.0245
R12326 avdd avdd.n447 0.0245
R12327 avdd.n443 avdd 0.0245
R12328 avdd avdd.n475 0.0245
R12329 avdd.n471 avdd 0.0245
R12330 avdd avdd.n503 0.0245
R12331 avdd.n499 avdd 0.0245
R12332 avdd avdd.n531 0.0245
R12333 avdd.n527 avdd 0.0245
R12334 avdd avdd.n559 0.0245
R12335 avdd.n555 avdd 0.0245
R12336 avdd avdd.n587 0.0245
R12337 avdd.n583 avdd 0.0245
R12338 avdd avdd.n615 0.0245
R12339 avdd.n611 avdd 0.0245
R12340 avdd avdd.n643 0.0245
R12341 avdd.n639 avdd 0.0245
R12342 avdd.n1194 avdd.n1171 0.0167304
R12343 avdd.n420 avdd.n408 0.016
R12344 avdd avdd.n1160 0.01225
R12345 avdd avdd.n64 0.012
R12346 avdd avdd.n56 0.012
R12347 avdd avdd.n48 0.012
R12348 avdd avdd.n40 0.012
R12349 avdd avdd.n32 0.012
R12350 avdd avdd.n24 0.012
R12351 avdd avdd.n16 0.012
R12352 avdd avdd.n8 0.012
R12353 avdd avdd.n0 0.012
R12354 avdd avdd.n401 0.012
R12355 avdd avdd.n393 0.012
R12356 avdd avdd.n385 0.012
R12357 avdd avdd.n377 0.012
R12358 avdd avdd.n369 0.012
R12359 avdd avdd.n361 0.012
R12360 avdd avdd.n353 0.012
R12361 avdd avdd.n345 0.012
R12362 avdd avdd.n337 0.012
R12363 avdd avdd.n78 0.009
R12364 avdd.n79 avdd 0.009
R12365 avdd.n91 avdd 0.009
R12366 avdd.n90 avdd 0.009
R12367 avdd.n89 avdd 0.009
R12368 avdd.n86 avdd 0.009
R12369 avdd.n110 avdd 0.009
R12370 avdd.n110 avdd 0.009
R12371 avdd.n109 avdd 0.009
R12372 avdd.n126 avdd 0.009
R12373 avdd.n125 avdd 0.009
R12374 avdd.n124 avdd 0.009
R12375 avdd.n118 avdd 0.009
R12376 avdd.n115 avdd 0.009
R12377 avdd.n138 avdd 0.009
R12378 avdd.n138 avdd 0.009
R12379 avdd.n137 avdd 0.009
R12380 avdd.n154 avdd 0.009
R12381 avdd.n153 avdd 0.009
R12382 avdd.n152 avdd 0.009
R12383 avdd.n146 avdd 0.009
R12384 avdd.n143 avdd 0.009
R12385 avdd.n166 avdd 0.009
R12386 avdd.n166 avdd 0.009
R12387 avdd.n165 avdd 0.009
R12388 avdd.n182 avdd 0.009
R12389 avdd.n181 avdd 0.009
R12390 avdd.n180 avdd 0.009
R12391 avdd.n174 avdd 0.009
R12392 avdd.n171 avdd 0.009
R12393 avdd.n194 avdd 0.009
R12394 avdd.n194 avdd 0.009
R12395 avdd.n193 avdd 0.009
R12396 avdd.n210 avdd 0.009
R12397 avdd.n209 avdd 0.009
R12398 avdd.n208 avdd 0.009
R12399 avdd.n202 avdd 0.009
R12400 avdd.n199 avdd 0.009
R12401 avdd.n222 avdd 0.009
R12402 avdd.n222 avdd 0.009
R12403 avdd.n221 avdd 0.009
R12404 avdd.n238 avdd 0.009
R12405 avdd.n237 avdd 0.009
R12406 avdd.n236 avdd 0.009
R12407 avdd.n230 avdd 0.009
R12408 avdd.n227 avdd 0.009
R12409 avdd.n250 avdd 0.009
R12410 avdd.n250 avdd 0.009
R12411 avdd.n249 avdd 0.009
R12412 avdd.n266 avdd 0.009
R12413 avdd.n265 avdd 0.009
R12414 avdd.n264 avdd 0.009
R12415 avdd.n258 avdd 0.009
R12416 avdd.n255 avdd 0.009
R12417 avdd.n278 avdd 0.009
R12418 avdd.n278 avdd 0.009
R12419 avdd.n277 avdd 0.009
R12420 avdd.n294 avdd 0.009
R12421 avdd.n293 avdd 0.009
R12422 avdd.n292 avdd 0.009
R12423 avdd.n286 avdd 0.009
R12424 avdd.n283 avdd 0.009
R12425 avdd.n306 avdd 0.009
R12426 avdd.n306 avdd 0.009
R12427 avdd.n305 avdd 0.009
R12428 avdd.n322 avdd 0.009
R12429 avdd.n321 avdd 0.009
R12430 avdd.n320 avdd 0.009
R12431 avdd.n314 avdd 0.009
R12432 avdd.n311 avdd 0.009
R12433 avdd.n334 avdd 0.009
R12434 avdd.n334 avdd 0.009
R12435 avdd.n333 avdd 0.009
R12436 avdd.n420 avdd 0.009
R12437 avdd.n419 avdd 0.009
R12438 avdd.n418 avdd 0.009
R12439 avdd.n415 avdd 0.009
R12440 avdd.n432 avdd 0.009
R12441 avdd.n432 avdd 0.009
R12442 avdd.n431 avdd 0.009
R12443 avdd.n448 avdd 0.009
R12444 avdd.n447 avdd 0.009
R12445 avdd.n446 avdd 0.009
R12446 avdd.n440 avdd 0.009
R12447 avdd.n437 avdd 0.009
R12448 avdd.n460 avdd 0.009
R12449 avdd.n460 avdd 0.009
R12450 avdd.n459 avdd 0.009
R12451 avdd.n476 avdd 0.009
R12452 avdd.n475 avdd 0.009
R12453 avdd.n474 avdd 0.009
R12454 avdd.n468 avdd 0.009
R12455 avdd.n465 avdd 0.009
R12456 avdd.n488 avdd 0.009
R12457 avdd.n488 avdd 0.009
R12458 avdd.n487 avdd 0.009
R12459 avdd.n504 avdd 0.009
R12460 avdd.n503 avdd 0.009
R12461 avdd.n502 avdd 0.009
R12462 avdd.n496 avdd 0.009
R12463 avdd.n493 avdd 0.009
R12464 avdd.n516 avdd 0.009
R12465 avdd.n516 avdd 0.009
R12466 avdd.n515 avdd 0.009
R12467 avdd.n532 avdd 0.009
R12468 avdd.n531 avdd 0.009
R12469 avdd.n530 avdd 0.009
R12470 avdd.n524 avdd 0.009
R12471 avdd.n521 avdd 0.009
R12472 avdd.n544 avdd 0.009
R12473 avdd.n544 avdd 0.009
R12474 avdd.n543 avdd 0.009
R12475 avdd.n560 avdd 0.009
R12476 avdd.n559 avdd 0.009
R12477 avdd.n558 avdd 0.009
R12478 avdd.n552 avdd 0.009
R12479 avdd.n549 avdd 0.009
R12480 avdd.n572 avdd 0.009
R12481 avdd.n572 avdd 0.009
R12482 avdd.n571 avdd 0.009
R12483 avdd.n588 avdd 0.009
R12484 avdd.n587 avdd 0.009
R12485 avdd.n586 avdd 0.009
R12486 avdd.n580 avdd 0.009
R12487 avdd.n577 avdd 0.009
R12488 avdd.n600 avdd 0.009
R12489 avdd.n600 avdd 0.009
R12490 avdd.n599 avdd 0.009
R12491 avdd.n616 avdd 0.009
R12492 avdd.n615 avdd 0.009
R12493 avdd.n614 avdd 0.009
R12494 avdd.n608 avdd 0.009
R12495 avdd.n605 avdd 0.009
R12496 avdd.n628 avdd 0.009
R12497 avdd.n628 avdd 0.009
R12498 avdd.n627 avdd 0.009
R12499 avdd.n644 avdd 0.009
R12500 avdd.n643 avdd 0.009
R12501 avdd.n642 avdd 0.009
R12502 avdd.n636 avdd 0.009
R12503 avdd.n633 avdd 0.009
R12504 avdd.n656 avdd 0.009
R12505 avdd.n656 avdd 0.009
R12506 avdd.n655 avdd 0.009
R12507 avdd avdd.n82 0.0085
R12508 avdd.n106 avdd.n105 0.0085
R12509 avdd.n134 avdd.n133 0.0085
R12510 avdd.n162 avdd.n161 0.0085
R12511 avdd.n190 avdd.n189 0.0085
R12512 avdd.n218 avdd.n217 0.0085
R12513 avdd.n246 avdd.n245 0.0085
R12514 avdd.n274 avdd.n273 0.0085
R12515 avdd.n302 avdd.n301 0.0085
R12516 avdd.n330 avdd.n329 0.0085
R12517 avdd.n428 avdd.n427 0.0085
R12518 avdd.n456 avdd.n455 0.0085
R12519 avdd.n484 avdd.n483 0.0085
R12520 avdd.n512 avdd.n511 0.0085
R12521 avdd.n540 avdd.n539 0.0085
R12522 avdd.n568 avdd.n567 0.0085
R12523 avdd.n596 avdd.n595 0.0085
R12524 avdd.n624 avdd.n623 0.0085
R12525 avdd.n652 avdd.n651 0.0085
R12526 avdd avdd.n89 0.0075
R12527 avdd.n118 avdd 0.0075
R12528 avdd.n146 avdd 0.0075
R12529 avdd.n174 avdd 0.0075
R12530 avdd.n202 avdd 0.0075
R12531 avdd.n230 avdd 0.0075
R12532 avdd.n258 avdd 0.0075
R12533 avdd.n286 avdd 0.0075
R12534 avdd.n314 avdd 0.0075
R12535 avdd avdd.n418 0.0075
R12536 avdd.n440 avdd 0.0075
R12537 avdd.n468 avdd 0.0075
R12538 avdd.n496 avdd 0.0075
R12539 avdd.n524 avdd 0.0075
R12540 avdd.n552 avdd 0.0075
R12541 avdd.n580 avdd 0.0075
R12542 avdd.n608 avdd 0.0075
R12543 avdd.n636 avdd 0.0075
R12544 avdd.n674 avdd.n662 0.00641216
R12545 avdd.n915 avdd.n914 0.00641216
R12546 avdd.n904 avdd.n903 0.00641216
R12547 avdd.n703 avdd.n700 0.00641216
R12548 avdd.n888 avdd.n706 0.00641216
R12549 avdd.n879 avdd.n878 0.00641216
R12550 avdd.n723 avdd.n720 0.00641216
R12551 avdd.n863 avdd.n726 0.00641216
R12552 avdd.n854 avdd.n853 0.00641216
R12553 avdd.n743 avdd.n740 0.00641216
R12554 avdd.n838 avdd.n746 0.00641216
R12555 avdd.n829 avdd.n828 0.00641216
R12556 avdd.n763 avdd.n760 0.00641216
R12557 avdd.n813 avdd.n766 0.00641216
R12558 avdd.n804 avdd.n803 0.00641216
R12559 avdd.n783 avdd.n780 0.00641216
R12560 avdd.n788 avdd.n787 0.00641216
R12561 avdd.n87 avdd 0.0055
R12562 avdd.n112 avdd.n64 0.0055
R12563 avdd.n120 avdd 0.0055
R12564 avdd.n140 avdd.n56 0.0055
R12565 avdd.n148 avdd 0.0055
R12566 avdd.n168 avdd.n48 0.0055
R12567 avdd.n176 avdd 0.0055
R12568 avdd.n196 avdd.n40 0.0055
R12569 avdd.n204 avdd 0.0055
R12570 avdd.n224 avdd.n32 0.0055
R12571 avdd.n232 avdd 0.0055
R12572 avdd.n252 avdd.n24 0.0055
R12573 avdd.n260 avdd 0.0055
R12574 avdd.n280 avdd.n16 0.0055
R12575 avdd.n288 avdd 0.0055
R12576 avdd.n308 avdd.n8 0.0055
R12577 avdd.n316 avdd 0.0055
R12578 avdd.n336 avdd.n0 0.0055
R12579 avdd.n416 avdd 0.0055
R12580 avdd.n434 avdd.n401 0.0055
R12581 avdd.n442 avdd 0.0055
R12582 avdd.n462 avdd.n393 0.0055
R12583 avdd.n470 avdd 0.0055
R12584 avdd.n490 avdd.n385 0.0055
R12585 avdd.n498 avdd 0.0055
R12586 avdd.n518 avdd.n377 0.0055
R12587 avdd.n526 avdd 0.0055
R12588 avdd.n546 avdd.n369 0.0055
R12589 avdd.n554 avdd 0.0055
R12590 avdd.n574 avdd.n361 0.0055
R12591 avdd.n582 avdd 0.0055
R12592 avdd.n602 avdd.n353 0.0055
R12593 avdd.n610 avdd 0.0055
R12594 avdd.n630 avdd.n345 0.0055
R12595 avdd.n638 avdd 0.0055
R12596 avdd.n658 avdd.n337 0.0055
R12597 avdd.n87 avdd.n85 0.004
R12598 avdd avdd.n112 0.004
R12599 avdd.n121 avdd.n120 0.004
R12600 avdd avdd.n140 0.004
R12601 avdd.n149 avdd.n148 0.004
R12602 avdd avdd.n168 0.004
R12603 avdd.n177 avdd.n176 0.004
R12604 avdd avdd.n196 0.004
R12605 avdd.n205 avdd.n204 0.004
R12606 avdd avdd.n224 0.004
R12607 avdd.n233 avdd.n232 0.004
R12608 avdd avdd.n252 0.004
R12609 avdd.n261 avdd.n260 0.004
R12610 avdd avdd.n280 0.004
R12611 avdd.n289 avdd.n288 0.004
R12612 avdd avdd.n308 0.004
R12613 avdd.n317 avdd.n316 0.004
R12614 avdd avdd.n336 0.004
R12615 avdd.n416 avdd.n414 0.004
R12616 avdd avdd.n434 0.004
R12617 avdd.n443 avdd.n442 0.004
R12618 avdd avdd.n462 0.004
R12619 avdd.n471 avdd.n470 0.004
R12620 avdd avdd.n490 0.004
R12621 avdd.n499 avdd.n498 0.004
R12622 avdd avdd.n518 0.004
R12623 avdd.n527 avdd.n526 0.004
R12624 avdd avdd.n546 0.004
R12625 avdd.n555 avdd.n554 0.004
R12626 avdd avdd.n574 0.004
R12627 avdd.n583 avdd.n582 0.004
R12628 avdd avdd.n602 0.004
R12629 avdd.n611 avdd.n610 0.004
R12630 avdd avdd.n630 0.004
R12631 avdd.n639 avdd.n638 0.004
R12632 avdd avdd.n658 0.004
R12633 avdd.n79 avdd 0.0035
R12634 avdd avdd.n109 0.003
R12635 avdd avdd.n137 0.003
R12636 avdd avdd.n165 0.003
R12637 avdd avdd.n193 0.003
R12638 avdd avdd.n221 0.003
R12639 avdd avdd.n249 0.003
R12640 avdd avdd.n277 0.003
R12641 avdd avdd.n305 0.003
R12642 avdd avdd.n333 0.003
R12643 avdd avdd.n431 0.003
R12644 avdd avdd.n459 0.003
R12645 avdd avdd.n487 0.003
R12646 avdd avdd.n515 0.003
R12647 avdd avdd.n543 0.003
R12648 avdd avdd.n571 0.003
R12649 avdd avdd.n599 0.003
R12650 avdd avdd.n627 0.003
R12651 avdd avdd.n655 0.003
R12652 avdd.n82 avdd.n81 0.001
R12653 avdd.n105 avdd 0.001
R12654 avdd.n133 avdd 0.001
R12655 avdd.n161 avdd 0.001
R12656 avdd.n189 avdd 0.001
R12657 avdd.n217 avdd 0.001
R12658 avdd.n245 avdd 0.001
R12659 avdd.n273 avdd 0.001
R12660 avdd.n301 avdd 0.001
R12661 avdd.n329 avdd 0.001
R12662 avdd.n427 avdd 0.001
R12663 avdd.n455 avdd 0.001
R12664 avdd.n483 avdd 0.001
R12665 avdd.n511 avdd 0.001
R12666 avdd.n539 avdd 0.001
R12667 avdd.n567 avdd 0.001
R12668 avdd.n595 avdd 0.001
R12669 avdd.n623 avdd 0.001
R12670 avdd.n651 avdd 0.001
R12671 otrip_decoded[0].n0 otrip_decoded[0].t1 186.374
R12672 otrip_decoded[0].n0 otrip_decoded[0].t0 170.308
R12673 otrip_decoded[0] otrip_decoded[0].n1 154.56
R12674 otrip_decoded[0].n2 otrip_decoded[0].n1 153.462
R12675 otrip_decoded[0].n1 otrip_decoded[0].n0 101.513
R12676 otrip_decoded[0].n3 otrip_decoded[0] 11.8005
R12677 otrip_decoded[0].n3 otrip_decoded[0].n2 4.96991
R12678 otrip_decoded[0].n2 otrip_decoded[0] 3.46403
R12679 otrip_decoded[0] otrip_decoded[0].n3 2.71109
R12680 rstring_mux_0.vtrip9.n2 rstring_mux_0.vtrip9.n0 50.7022
R12681 rstring_mux_0.vtrip9.n2 rstring_mux_0.vtrip9.n1 13.8791
R12682 rstring_mux_0.vtrip9.t2 rstring_mux_0.vtrip9.n3 10.5857
R12683 rstring_mux_0.vtrip9.n3 rstring_mux_0.vtrip9.t5 10.5847
R12684 rstring_mux_0.vtrip9.n3 rstring_mux_0.vtrip9.n2 8.35755
R12685 rstring_mux_0.vtrip9.n0 rstring_mux_0.vtrip9.t4 5.5395
R12686 rstring_mux_0.vtrip9.n0 rstring_mux_0.vtrip9.t3 5.5395
R12687 rstring_mux_0.vtrip9.n1 rstring_mux_0.vtrip9.t0 3.3065
R12688 rstring_mux_0.vtrip9.n1 rstring_mux_0.vtrip9.t1 3.3065
R12689 rstring_mux_0.vtrip8.n2 rstring_mux_0.vtrip8.n0 50.7022
R12690 rstring_mux_0.vtrip8.n3 rstring_mux_0.vtrip8.n2 16.7526
R12691 rstring_mux_0.vtrip8.n2 rstring_mux_0.vtrip8.n1 13.8791
R12692 rstring_mux_0.vtrip8.n3 rstring_mux_0.vtrip8.t3 10.6303
R12693 rstring_mux_0.vtrip8.n0 rstring_mux_0.vtrip8.t5 5.5395
R12694 rstring_mux_0.vtrip8.n0 rstring_mux_0.vtrip8.t4 5.5395
R12695 rstring_mux_0.vtrip8.n1 rstring_mux_0.vtrip8.t0 3.3065
R12696 rstring_mux_0.vtrip8.n1 rstring_mux_0.vtrip8.t1 3.3065
R12697 rstring_mux_0.vtrip8.t2 rstring_mux_0.vtrip8.n3 0.825482
R12698 schmitt_trigger_0.out.n8 schmitt_trigger_0.out.t8 248.236
R12699 schmitt_trigger_0.out.n6 schmitt_trigger_0.out.t6 240.778
R12700 schmitt_trigger_0.out.n7 schmitt_trigger_0.out.t15 240.613
R12701 schmitt_trigger_0.out.n6 schmitt_trigger_0.out.t12 240.349
R12702 schmitt_trigger_0.out.n5 schmitt_trigger_0.out.t0 236.369
R12703 schmitt_trigger_0.out.n0 schmitt_trigger_0.out.t5 212.081
R12704 schmitt_trigger_0.out.n2 schmitt_trigger_0.out.t4 212.081
R12705 schmitt_trigger_0.out.n15 schmitt_trigger_0.out.t7 212.081
R12706 schmitt_trigger_0.out.n3 schmitt_trigger_0.out.t14 212.081
R12707 schmitt_trigger_0.out.n5 schmitt_trigger_0.out.n4 207.585
R12708 schmitt_trigger_0.out.n12 schmitt_trigger_0.out.n3 188.516
R12709 sky130_fd_sc_hd__inv_4_0.A schmitt_trigger_0.out.n1 154.304
R12710 schmitt_trigger_0.out.n14 schmitt_trigger_0.out.n13 152
R12711 schmitt_trigger_0.out.n17 schmitt_trigger_0.out.n16 152
R12712 schmitt_trigger_0.out.n0 schmitt_trigger_0.out.t11 139.78
R12713 schmitt_trigger_0.out.n2 schmitt_trigger_0.out.t10 139.78
R12714 schmitt_trigger_0.out.n15 schmitt_trigger_0.out.t13 139.78
R12715 schmitt_trigger_0.out.n3 schmitt_trigger_0.out.t9 139.78
R12716 schmitt_trigger_0.out.n10 schmitt_trigger_0.out.t3 91.727
R12717 schmitt_trigger_0.out.n1 schmitt_trigger_0.out.n0 30.6732
R12718 schmitt_trigger_0.out.n2 schmitt_trigger_0.out.n1 30.6732
R12719 schmitt_trigger_0.out.n16 schmitt_trigger_0.out.n2 30.6732
R12720 schmitt_trigger_0.out.n16 schmitt_trigger_0.out.n15 30.6732
R12721 schmitt_trigger_0.out.n15 schmitt_trigger_0.out.n14 30.6732
R12722 schmitt_trigger_0.out.n14 schmitt_trigger_0.out.n3 30.6732
R12723 schmitt_trigger_0.out.n4 schmitt_trigger_0.out.t1 28.5655
R12724 schmitt_trigger_0.out.n4 schmitt_trigger_0.out.t2 28.5655
R12725 schmitt_trigger_0.out.n11 schmitt_trigger_0.out.n10 20.1312
R12726 sky130_fd_sc_hd__inv_4_0.A schmitt_trigger_0.out.n17 19.2005
R12727 sky130_fd_sc_hd__inv_4_0.A schmitt_trigger_0.out.n12 17.1525
R12728 schmitt_trigger_0.out.n11 sky130_fd_sc_hd__inv_4_0.A 12.8005
R12729 schmitt_trigger_0.out.n9 schmitt_trigger_0.out.n5 8.66251
R12730 schmitt_trigger_0.out.n13 sky130_fd_sc_hd__inv_4_0.A 6.4005
R12731 schmitt_trigger_0.out.n12 sky130_fd_sc_hd__inv_4_0.A 6.4005
R12732 schmitt_trigger_0.out.n8 schmitt_trigger_0.out.n7 4.94425
R12733 schmitt_trigger_0.out.n17 sky130_fd_sc_hd__inv_4_0.A 4.3525
R12734 schmitt_trigger_0.out.n13 schmitt_trigger_0.out.n11 4.3525
R12735 schmitt_trigger_0.out.n9 schmitt_trigger_0.out.n8 4.05633
R12736 schmitt_trigger_0.out.n10 schmitt_trigger_0.out.n9 0.230017
R12737 schmitt_trigger_0.out.n7 schmitt_trigger_0.out.n6 0.117348
R12738 dvdd.n186 dvdd.n183 15967.3
R12739 dvdd.n187 dvdd.n186 15967.3
R12740 dvdd.n188 dvdd.n183 15967.3
R12741 dvdd.n188 dvdd.n187 15967.3
R12742 dvdd.n185 dvdd.n181 8190.81
R12743 dvdd.n185 dvdd.n182 8190.81
R12744 dvdd.n189 dvdd.n181 8190.81
R12745 dvdd.n189 dvdd.n182 8190.81
R12746 dvdd.n117 dvdd.n116 4782.35
R12747 dvdd.n118 dvdd.n116 4782.35
R12748 dvdd.n117 dvdd.n101 4782.35
R12749 dvdd.n118 dvdd.n101 4782.35
R12750 dvdd.n184 dvdd.n179 1909.08
R12751 dvdd.n184 dvdd.n180 1909.08
R12752 dvdd.n190 dvdd.n180 1909.08
R12753 dvdd.n191 dvdd.n190 1723.48
R12754 dvdd.n170 dvdd.t71 871.962
R12755 dvdd.n119 dvdd.n115 510.118
R12756 dvdd.n120 dvdd.n119 510.118
R12757 dvdd.n120 dvdd.n100 510.118
R12758 dvdd.n115 dvdd.n100 510.118
R12759 dvdd.t102 dvdd.n117 369.05
R12760 dvdd.n118 dvdd.t22 369.05
R12761 dvdd.n137 dvdd.t43 348.805
R12762 dvdd dvdd.t70 336.933
R12763 dvdd.n175 dvdd.n124 320.976
R12764 dvdd.n164 dvdd.n128 320.976
R12765 dvdd.n130 dvdd.n129 320.976
R12766 dvdd.n156 dvdd.n132 320.976
R12767 dvdd.n150 dvdd.n149 320.976
R12768 dvdd.n147 dvdd.n135 320.976
R12769 dvdd.n141 dvdd.n140 320.976
R12770 dvdd.n139 dvdd.n138 320.976
R12771 dvdd.n300 dvdd.n194 307.762
R12772 dvdd.n296 dvdd.n201 307.762
R12773 dvdd.n292 dvdd.n208 307.762
R12774 dvdd.n288 dvdd.n215 307.762
R12775 dvdd.n284 dvdd.n222 307.762
R12776 dvdd.n280 dvdd.n229 307.762
R12777 dvdd.n276 dvdd.n236 307.762
R12778 dvdd.n272 dvdd.n243 307.762
R12779 dvdd.n268 dvdd.n250 307.762
R12780 dvdd.n96 dvdd.n0 307.762
R12781 dvdd.n92 dvdd.n7 307.762
R12782 dvdd.n88 dvdd.n14 307.762
R12783 dvdd.n84 dvdd.n21 307.762
R12784 dvdd.n80 dvdd.n28 307.762
R12785 dvdd.n76 dvdd.n35 307.762
R12786 dvdd.n72 dvdd.n42 307.762
R12787 dvdd.n68 dvdd.n49 307.762
R12788 dvdd.n64 dvdd.n56 307.762
R12789 dvdd.t104 dvdd.t102 264.262
R12790 dvdd.t106 dvdd.t104 264.262
R12791 dvdd.t121 dvdd.t106 264.262
R12792 dvdd.t68 dvdd.t121 264.262
R12793 dvdd.t64 dvdd.t68 264.262
R12794 dvdd.t60 dvdd.t64 264.262
R12795 dvdd.t16 dvdd.t60 264.262
R12796 dvdd.t18 dvdd.t16 264.262
R12797 dvdd.t24 dvdd.t18 264.262
R12798 dvdd.t14 dvdd.t24 264.262
R12799 dvdd.t20 dvdd.t14 264.262
R12800 dvdd.t22 dvdd.t20 264.262
R12801 dvdd.n126 dvdd.t55 250.785
R12802 dvdd.n262 dvdd.t113 246.106
R12803 dvdd.n177 dvdd.t63 244.737
R12804 dvdd.n99 dvdd.t120 240.488
R12805 dvdd.n98 dvdd.t23 228.669
R12806 dvdd.t56 dvdd.t42 212.8
R12807 dvdd.t36 dvdd.t56 212.8
R12808 dvdd.t48 dvdd.t36 212.8
R12809 dvdd.t40 dvdd.t48 212.8
R12810 dvdd.t28 dvdd.t40 212.8
R12811 dvdd.t30 dvdd.t28 212.8
R12812 dvdd.t52 dvdd.t30 212.8
R12813 dvdd.t58 dvdd.t52 212.8
R12814 dvdd.t44 dvdd.t58 212.8
R12815 dvdd.t34 dvdd.t44 212.8
R12816 dvdd.t46 dvdd.t38 212.8
R12817 dvdd.t38 dvdd.t50 212.8
R12818 dvdd.t50 dvdd.t32 212.8
R12819 dvdd.t32 dvdd.t54 212.8
R12820 dvdd.t70 dvdd.t72 212.8
R12821 dvdd.t72 dvdd.t66 212.8
R12822 dvdd.t66 dvdd.t62 212.8
R12823 dvdd.n264 dvdd.n257 205.5
R12824 dvdd.n111 dvdd.n110 200.105
R12825 dvdd.n112 dvdd.n109 200.105
R12826 dvdd.n113 dvdd.n108 200.105
R12827 dvdd.n107 dvdd.n102 200.105
R12828 dvdd.n106 dvdd.n103 200.105
R12829 dvdd.n105 dvdd.n104 200.105
R12830 dvdd.t54 dvdd 197.601
R12831 dvdd.t62 dvdd 190
R12832 dvdd.n198 dvdd.n195 185
R12833 dvdd.n199 dvdd.n198 185
R12834 dvdd.n205 dvdd.n202 185
R12835 dvdd.n206 dvdd.n205 185
R12836 dvdd.n212 dvdd.n209 185
R12837 dvdd.n213 dvdd.n212 185
R12838 dvdd.n219 dvdd.n216 185
R12839 dvdd.n220 dvdd.n219 185
R12840 dvdd.n226 dvdd.n223 185
R12841 dvdd.n227 dvdd.n226 185
R12842 dvdd.n233 dvdd.n230 185
R12843 dvdd.n234 dvdd.n233 185
R12844 dvdd.n240 dvdd.n237 185
R12845 dvdd.n241 dvdd.n240 185
R12846 dvdd.n247 dvdd.n244 185
R12847 dvdd.n248 dvdd.n247 185
R12848 dvdd.n254 dvdd.n251 185
R12849 dvdd.n255 dvdd.n254 185
R12850 dvdd.n4 dvdd.n1 185
R12851 dvdd.n5 dvdd.n4 185
R12852 dvdd.n11 dvdd.n8 185
R12853 dvdd.n12 dvdd.n11 185
R12854 dvdd.n18 dvdd.n15 185
R12855 dvdd.n19 dvdd.n18 185
R12856 dvdd.n25 dvdd.n22 185
R12857 dvdd.n26 dvdd.n25 185
R12858 dvdd.n32 dvdd.n29 185
R12859 dvdd.n33 dvdd.n32 185
R12860 dvdd.n39 dvdd.n36 185
R12861 dvdd.n40 dvdd.n39 185
R12862 dvdd.n46 dvdd.n43 185
R12863 dvdd.n47 dvdd.n46 185
R12864 dvdd.n53 dvdd.n50 185
R12865 dvdd.n54 dvdd.n53 185
R12866 dvdd.n60 dvdd.n57 185
R12867 dvdd.n61 dvdd.n60 185
R12868 dvdd.n191 dvdd.n179 166.776
R12869 dvdd.n261 dvdd.t112 157.446
R12870 dvdd.n158 dvdd.t46 141.868
R12871 dvdd.t10 dvdd.n197 129.546
R12872 dvdd.t134 dvdd.n204 129.546
R12873 dvdd.t26 dvdd.n211 129.546
R12874 dvdd.t142 dvdd.n218 129.546
R12875 dvdd.t76 dvdd.n225 129.546
R12876 dvdd.t82 dvdd.n232 129.546
R12877 dvdd.t140 dvdd.n239 129.546
R12878 dvdd.t8 dvdd.n246 129.546
R12879 dvdd.t6 dvdd.n253 129.546
R12880 dvdd.t84 dvdd.n3 129.546
R12881 dvdd.t136 dvdd.n10 129.546
R12882 dvdd.t78 dvdd.n17 129.546
R12883 dvdd.t108 dvdd.n24 129.546
R12884 dvdd.t74 dvdd.n31 129.546
R12885 dvdd.t90 dvdd.n38 129.546
R12886 dvdd.t110 dvdd.n45 129.546
R12887 dvdd.t118 dvdd.n52 129.546
R12888 dvdd.t88 dvdd.n59 129.546
R12889 dvdd.t131 dvdd.n258 127.638
R12890 dvdd.n200 dvdd.n195 101.644
R12891 dvdd.n207 dvdd.n202 101.644
R12892 dvdd.n214 dvdd.n209 101.644
R12893 dvdd.n221 dvdd.n216 101.644
R12894 dvdd.n228 dvdd.n223 101.644
R12895 dvdd.n235 dvdd.n230 101.644
R12896 dvdd.n242 dvdd.n237 101.644
R12897 dvdd.n249 dvdd.n244 101.644
R12898 dvdd.n256 dvdd.n251 101.644
R12899 dvdd.n6 dvdd.n1 101.644
R12900 dvdd.n13 dvdd.n8 101.644
R12901 dvdd.n20 dvdd.n15 101.644
R12902 dvdd.n27 dvdd.n22 101.644
R12903 dvdd.n34 dvdd.n29 101.644
R12904 dvdd.n41 dvdd.n36 101.644
R12905 dvdd.n48 dvdd.n43 101.644
R12906 dvdd.n55 dvdd.n50 101.644
R12907 dvdd.n62 dvdd.n57 101.644
R12908 dvdd.n263 dvdd.n258 95.8438
R12909 dvdd.n260 dvdd.n259 92.5005
R12910 dvdd.n200 dvdd.n199 92.5005
R12911 dvdd.n207 dvdd.n206 92.5005
R12912 dvdd.n214 dvdd.n213 92.5005
R12913 dvdd.n221 dvdd.n220 92.5005
R12914 dvdd.n228 dvdd.n227 92.5005
R12915 dvdd.n235 dvdd.n234 92.5005
R12916 dvdd.n242 dvdd.n241 92.5005
R12917 dvdd.n249 dvdd.n248 92.5005
R12918 dvdd.n256 dvdd.n255 92.5005
R12919 dvdd.n6 dvdd.n5 92.5005
R12920 dvdd.n13 dvdd.n12 92.5005
R12921 dvdd.n20 dvdd.n19 92.5005
R12922 dvdd.n27 dvdd.n26 92.5005
R12923 dvdd.n34 dvdd.n33 92.5005
R12924 dvdd.n41 dvdd.n40 92.5005
R12925 dvdd.n48 dvdd.n47 92.5005
R12926 dvdd.n55 dvdd.n54 92.5005
R12927 dvdd.n62 dvdd.n61 92.5005
R12928 dvdd.n260 dvdd.n258 82.3534
R12929 dvdd.n197 dvdd.n196 77.057
R12930 dvdd.n204 dvdd.n203 77.057
R12931 dvdd.n211 dvdd.n210 77.057
R12932 dvdd.n218 dvdd.n217 77.057
R12933 dvdd.n225 dvdd.n224 77.057
R12934 dvdd.n232 dvdd.n231 77.057
R12935 dvdd.n239 dvdd.n238 77.057
R12936 dvdd.n246 dvdd.n245 77.057
R12937 dvdd.n253 dvdd.n252 77.057
R12938 dvdd.n3 dvdd.n2 77.057
R12939 dvdd.n10 dvdd.n9 77.057
R12940 dvdd.n17 dvdd.n16 77.057
R12941 dvdd.n24 dvdd.n23 77.057
R12942 dvdd.n31 dvdd.n30 77.057
R12943 dvdd.n38 dvdd.n37 77.057
R12944 dvdd.n45 dvdd.n44 77.057
R12945 dvdd.n52 dvdd.n51 77.057
R12946 dvdd.n59 dvdd.n58 77.057
R12947 dvdd.n158 dvdd.t34 70.9338
R12948 dvdd.n198 dvdd.t10 67.8576
R12949 dvdd.n205 dvdd.t134 67.8576
R12950 dvdd.n212 dvdd.t26 67.8576
R12951 dvdd.n219 dvdd.t142 67.8576
R12952 dvdd.n226 dvdd.t76 67.8576
R12953 dvdd.n233 dvdd.t82 67.8576
R12954 dvdd.n240 dvdd.t140 67.8576
R12955 dvdd.n247 dvdd.t8 67.8576
R12956 dvdd.n254 dvdd.t6 67.8576
R12957 dvdd.n4 dvdd.t84 67.8576
R12958 dvdd.n11 dvdd.t136 67.8576
R12959 dvdd.n18 dvdd.t78 67.8576
R12960 dvdd.n25 dvdd.t108 67.8576
R12961 dvdd.n32 dvdd.t74 67.8576
R12962 dvdd.n39 dvdd.t90 67.8576
R12963 dvdd.n46 dvdd.t110 67.8576
R12964 dvdd.n53 dvdd.t118 67.8576
R12965 dvdd.n60 dvdd.t88 67.8576
R12966 dvdd.n259 dvdd.t131 55.9594
R12967 dvdd.n259 dvdd.t112 55.9594
R12968 dvdd.n197 dvdd.t12 47.2949
R12969 dvdd.n204 dvdd.t127 47.2949
R12970 dvdd.n211 dvdd.t129 47.2949
R12971 dvdd.n218 dvdd.t114 47.2949
R12972 dvdd.n225 dvdd.t0 47.2949
R12973 dvdd.n232 dvdd.t86 47.2949
R12974 dvdd.n239 dvdd.t123 47.2949
R12975 dvdd.n246 dvdd.t98 47.2949
R12976 dvdd.n253 dvdd.t2 47.2949
R12977 dvdd.n3 dvdd.t4 47.2949
R12978 dvdd.n10 dvdd.t125 47.2949
R12979 dvdd.n17 dvdd.t138 47.2949
R12980 dvdd.n24 dvdd.t100 47.2949
R12981 dvdd.n31 dvdd.t94 47.2949
R12982 dvdd.n38 dvdd.t92 47.2949
R12983 dvdd.n45 dvdd.t116 47.2949
R12984 dvdd.n52 dvdd.t80 47.2949
R12985 dvdd.n59 dvdd.t96 47.2949
R12986 dvdd.n119 dvdd.n118 46.2505
R12987 dvdd.n117 dvdd.n100 46.2505
R12988 dvdd.n262 dvdd.n261 33.4807
R12989 dvdd.n194 dvdd.t11 32.8338
R12990 dvdd.n194 dvdd.t13 32.8338
R12991 dvdd.n201 dvdd.t135 32.8338
R12992 dvdd.n201 dvdd.t128 32.8338
R12993 dvdd.n208 dvdd.t27 32.8338
R12994 dvdd.n208 dvdd.t130 32.8338
R12995 dvdd.n215 dvdd.t143 32.8338
R12996 dvdd.n215 dvdd.t115 32.8338
R12997 dvdd.n222 dvdd.t77 32.8338
R12998 dvdd.n222 dvdd.t1 32.8338
R12999 dvdd.n229 dvdd.t83 32.8338
R13000 dvdd.n229 dvdd.t87 32.8338
R13001 dvdd.n236 dvdd.t141 32.8338
R13002 dvdd.n236 dvdd.t124 32.8338
R13003 dvdd.n243 dvdd.t9 32.8338
R13004 dvdd.n243 dvdd.t99 32.8338
R13005 dvdd.n250 dvdd.t7 32.8338
R13006 dvdd.n250 dvdd.t3 32.8338
R13007 dvdd.n0 dvdd.t85 32.8338
R13008 dvdd.n0 dvdd.t5 32.8338
R13009 dvdd.n7 dvdd.t137 32.8338
R13010 dvdd.n7 dvdd.t126 32.8338
R13011 dvdd.n14 dvdd.t79 32.8338
R13012 dvdd.n14 dvdd.t139 32.8338
R13013 dvdd.n21 dvdd.t109 32.8338
R13014 dvdd.n21 dvdd.t101 32.8338
R13015 dvdd.n28 dvdd.t75 32.8338
R13016 dvdd.n28 dvdd.t95 32.8338
R13017 dvdd.n35 dvdd.t91 32.8338
R13018 dvdd.n35 dvdd.t93 32.8338
R13019 dvdd.n42 dvdd.t111 32.8338
R13020 dvdd.n42 dvdd.t117 32.8338
R13021 dvdd.n49 dvdd.t119 32.8338
R13022 dvdd.n49 dvdd.t81 32.8338
R13023 dvdd.n56 dvdd.t89 32.8338
R13024 dvdd.n56 dvdd.t97 32.8338
R13025 dvdd.n199 dvdd.n196 30.8889
R13026 dvdd.n196 dvdd.n195 30.8889
R13027 dvdd.n206 dvdd.n203 30.8889
R13028 dvdd.n203 dvdd.n202 30.8889
R13029 dvdd.n213 dvdd.n210 30.8889
R13030 dvdd.n210 dvdd.n209 30.8889
R13031 dvdd.n220 dvdd.n217 30.8889
R13032 dvdd.n217 dvdd.n216 30.8889
R13033 dvdd.n227 dvdd.n224 30.8889
R13034 dvdd.n224 dvdd.n223 30.8889
R13035 dvdd.n234 dvdd.n231 30.8889
R13036 dvdd.n231 dvdd.n230 30.8889
R13037 dvdd.n241 dvdd.n238 30.8889
R13038 dvdd.n238 dvdd.n237 30.8889
R13039 dvdd.n248 dvdd.n245 30.8889
R13040 dvdd.n245 dvdd.n244 30.8889
R13041 dvdd.n255 dvdd.n252 30.8889
R13042 dvdd.n252 dvdd.n251 30.8889
R13043 dvdd.n5 dvdd.n2 30.8889
R13044 dvdd.n2 dvdd.n1 30.8889
R13045 dvdd.n12 dvdd.n9 30.8889
R13046 dvdd.n9 dvdd.n8 30.8889
R13047 dvdd.n19 dvdd.n16 30.8889
R13048 dvdd.n16 dvdd.n15 30.8889
R13049 dvdd.n26 dvdd.n23 30.8889
R13050 dvdd.n23 dvdd.n22 30.8889
R13051 dvdd.n33 dvdd.n30 30.8889
R13052 dvdd.n30 dvdd.n29 30.8889
R13053 dvdd.n40 dvdd.n37 30.8889
R13054 dvdd.n37 dvdd.n36 30.8889
R13055 dvdd.n47 dvdd.n44 30.8889
R13056 dvdd.n44 dvdd.n43 30.8889
R13057 dvdd.n54 dvdd.n51 30.8889
R13058 dvdd.n51 dvdd.n50 30.8889
R13059 dvdd.n61 dvdd.n58 30.8889
R13060 dvdd.n58 dvdd.n57 30.8889
R13061 dvdd.n110 dvdd.t15 28.5655
R13062 dvdd.n110 dvdd.t21 28.5655
R13063 dvdd.n109 dvdd.t19 28.5655
R13064 dvdd.n109 dvdd.t25 28.5655
R13065 dvdd.n108 dvdd.t61 28.5655
R13066 dvdd.n108 dvdd.t17 28.5655
R13067 dvdd.n102 dvdd.t69 28.5655
R13068 dvdd.n102 dvdd.t65 28.5655
R13069 dvdd.n103 dvdd.t107 28.5655
R13070 dvdd.n103 dvdd.t122 28.5655
R13071 dvdd.n104 dvdd.t103 28.5655
R13072 dvdd.n104 dvdd.t105 28.5655
R13073 dvdd.n261 dvdd.n260 27.7986
R13074 dvdd.n124 dvdd.t73 26.5955
R13075 dvdd.n124 dvdd.t67 26.5955
R13076 dvdd.n128 dvdd.t51 26.5955
R13077 dvdd.n128 dvdd.t33 26.5955
R13078 dvdd.n129 dvdd.t47 26.5955
R13079 dvdd.n129 dvdd.t39 26.5955
R13080 dvdd.n132 dvdd.t45 26.5955
R13081 dvdd.n132 dvdd.t35 26.5955
R13082 dvdd.n149 dvdd.t53 26.5955
R13083 dvdd.n149 dvdd.t59 26.5955
R13084 dvdd.n135 dvdd.t29 26.5955
R13085 dvdd.n135 dvdd.t31 26.5955
R13086 dvdd.n140 dvdd.t49 26.5955
R13087 dvdd.n140 dvdd.t41 26.5955
R13088 dvdd.n138 dvdd.t57 26.5955
R13089 dvdd.n138 dvdd.t37 26.5955
R13090 dvdd.n257 dvdd.t132 24.6255
R13091 dvdd.n257 dvdd.t133 24.6255
R13092 dvdd.n63 dvdd 22.5644
R13093 dvdd.n299 dvdd.n298 22.5272
R13094 dvdd.n295 dvdd.n294 22.5272
R13095 dvdd.n291 dvdd.n290 22.5272
R13096 dvdd.n287 dvdd.n286 22.5272
R13097 dvdd.n283 dvdd.n282 22.5272
R13098 dvdd.n279 dvdd.n278 22.5272
R13099 dvdd.n275 dvdd.n274 22.5272
R13100 dvdd.n271 dvdd.n270 22.5272
R13101 dvdd.n267 dvdd.n266 22.5272
R13102 dvdd.n95 dvdd.n94 22.5272
R13103 dvdd.n91 dvdd.n90 22.5272
R13104 dvdd.n87 dvdd.n86 22.5272
R13105 dvdd.n83 dvdd.n82 22.5272
R13106 dvdd.n79 dvdd.n78 22.5272
R13107 dvdd.n75 dvdd.n74 22.5272
R13108 dvdd.n71 dvdd.n70 22.5272
R13109 dvdd.n67 dvdd.n66 22.5272
R13110 dvdd.n300 dvdd.n299 17.4938
R13111 dvdd.n296 dvdd.n295 17.4938
R13112 dvdd.n292 dvdd.n291 17.4938
R13113 dvdd.n288 dvdd.n287 17.4938
R13114 dvdd.n284 dvdd.n283 17.4938
R13115 dvdd.n280 dvdd.n279 17.4938
R13116 dvdd.n276 dvdd.n275 17.4938
R13117 dvdd.n272 dvdd.n271 17.4938
R13118 dvdd.n268 dvdd.n267 17.4938
R13119 dvdd.n96 dvdd.n95 17.4938
R13120 dvdd.n92 dvdd.n91 17.4938
R13121 dvdd.n88 dvdd.n87 17.4938
R13122 dvdd.n84 dvdd.n83 17.4938
R13123 dvdd.n80 dvdd.n79 17.4938
R13124 dvdd.n76 dvdd.n75 17.4938
R13125 dvdd.n72 dvdd.n71 17.4938
R13126 dvdd.n68 dvdd.n67 17.4938
R13127 dvdd.n64 dvdd.n63 17.4938
R13128 dvdd.n146 dvdd.n136 16.132
R13129 dvdd.n151 dvdd.n148 16.132
R13130 dvdd.n155 dvdd.n133 16.132
R13131 dvdd.n166 dvdd.n165 16.132
R13132 dvdd.n171 dvdd.n169 16.132
R13133 dvdd.n175 dvdd.n125 16.132
R13134 dvdd.n176 dvdd.n175 16.132
R13135 dvdd.n142 dvdd.n139 15.9567
R13136 dvdd.n164 dvdd.n163 15.606
R13137 dvdd.n263 dvdd 15.5495
R13138 dvdd.n177 dvdd.n176 15.08
R13139 dvdd.n160 dvdd.n159 14.9046
R13140 dvdd.n159 dvdd.n158 14.2313
R13141 dvdd.n170 dvdd.n125 14.0279
R13142 dvdd.n163 dvdd.n130 13.8526
R13143 dvdd.n142 dvdd.n141 13.5019
R13144 dvdd.n166 dvdd.n126 13.5019
R13145 dvdd.n157 dvdd.n156 11.0471
R13146 dvdd.n302 dvdd.n193 10.8092
R13147 dvdd.n147 dvdd.n146 10.6964
R13148 dvdd.n178 dvdd.n177 10.3526
R13149 dvdd.n265 dvdd.n264 10.0534
R13150 dvdd.n192 dvdd.n191 9.45415
R13151 dvdd.n143 dvdd.n142 9.3005
R13152 dvdd.n144 dvdd.n136 9.3005
R13153 dvdd.n146 dvdd.n145 9.3005
R13154 dvdd.n148 dvdd.n134 9.3005
R13155 dvdd.n152 dvdd.n151 9.3005
R13156 dvdd.n153 dvdd.n133 9.3005
R13157 dvdd.n155 dvdd.n154 9.3005
R13158 dvdd.n157 dvdd.n131 9.3005
R13159 dvdd.n161 dvdd.n160 9.3005
R13160 dvdd.n163 dvdd.n162 9.3005
R13161 dvdd.n165 dvdd.n127 9.3005
R13162 dvdd.n167 dvdd.n166 9.3005
R13163 dvdd.n169 dvdd.n168 9.3005
R13164 dvdd.n172 dvdd.n171 9.3005
R13165 dvdd.n173 dvdd.n125 9.3005
R13166 dvdd.n175 dvdd.n174 9.3005
R13167 dvdd.n176 dvdd.n123 9.3005
R13168 dvdd.n269 dvdd.n268 9.3005
R13169 dvdd.n273 dvdd.n272 9.3005
R13170 dvdd.n277 dvdd.n276 9.3005
R13171 dvdd.n281 dvdd.n280 9.3005
R13172 dvdd.n285 dvdd.n284 9.3005
R13173 dvdd.n289 dvdd.n288 9.3005
R13174 dvdd.n293 dvdd.n292 9.3005
R13175 dvdd.n297 dvdd.n296 9.3005
R13176 dvdd.n301 dvdd.n300 9.3005
R13177 dvdd.n65 dvdd.n64 9.3005
R13178 dvdd.n69 dvdd.n68 9.3005
R13179 dvdd.n73 dvdd.n72 9.3005
R13180 dvdd.n77 dvdd.n76 9.3005
R13181 dvdd.n81 dvdd.n80 9.3005
R13182 dvdd.n85 dvdd.n84 9.3005
R13183 dvdd.n89 dvdd.n88 9.3005
R13184 dvdd.n93 dvdd.n92 9.3005
R13185 dvdd.n97 dvdd.n96 9.3005
R13186 dvdd.n150 dvdd.n133 8.2416
R13187 dvdd.n151 dvdd.n150 7.89091
R13188 dvdd.n264 dvdd.n263 6.58874
R13189 dvdd.n120 dvdd.n101 5.96824
R13190 dvdd.t60 dvdd.n101 5.96824
R13191 dvdd.n116 dvdd.n115 5.96824
R13192 dvdd.t60 dvdd.n116 5.96824
R13193 dvdd.n139 dvdd.n137 5.87299
R13194 dvdd.n148 dvdd.n147 5.43612
R13195 dvdd.n156 dvdd.n155 5.08543
R13196 dvdd.n303 dvdd 5.04667
R13197 dvdd.n193 dvdd.n192 4.5005
R13198 dvdd.n299 dvdd.n200 4.32258
R13199 dvdd.n295 dvdd.n207 4.32258
R13200 dvdd.n291 dvdd.n214 4.32258
R13201 dvdd.n287 dvdd.n221 4.32258
R13202 dvdd.n283 dvdd.n228 4.32258
R13203 dvdd.n279 dvdd.n235 4.32258
R13204 dvdd.n275 dvdd.n242 4.32258
R13205 dvdd.n271 dvdd.n249 4.32258
R13206 dvdd.n267 dvdd.n256 4.32258
R13207 dvdd.n95 dvdd.n6 4.32258
R13208 dvdd.n91 dvdd.n13 4.32258
R13209 dvdd.n87 dvdd.n20 4.32258
R13210 dvdd.n83 dvdd.n27 4.32258
R13211 dvdd.n79 dvdd.n34 4.32258
R13212 dvdd.n75 dvdd.n41 4.32258
R13213 dvdd.n71 dvdd.n48 4.32258
R13214 dvdd.n67 dvdd.n55 4.32258
R13215 dvdd.n63 dvdd.n62 4.32258
R13216 dvdd.n193 dvdd.n122 3.79251
R13217 dvdd.n302 dvdd 3.73954
R13218 dvdd dvdd.n303 3.73954
R13219 dvdd.n185 dvdd.n184 3.7005
R13220 dvdd.n186 dvdd.n185 3.7005
R13221 dvdd.n190 dvdd.n189 3.7005
R13222 dvdd.n189 dvdd.n188 3.7005
R13223 dvdd.n122 dvdd.n121 3.36211
R13224 dvdd.n263 dvdd.n262 3.34378
R13225 dvdd.n266 dvdd 2.9391
R13226 dvdd.n270 dvdd 2.9391
R13227 dvdd.n274 dvdd 2.9391
R13228 dvdd.n278 dvdd 2.9391
R13229 dvdd.n282 dvdd 2.9391
R13230 dvdd.n286 dvdd 2.9391
R13231 dvdd.n290 dvdd 2.9391
R13232 dvdd.n294 dvdd 2.9391
R13233 dvdd.n298 dvdd 2.9391
R13234 dvdd.n66 dvdd 2.9391
R13235 dvdd.n70 dvdd 2.9391
R13236 dvdd.n74 dvdd 2.9391
R13237 dvdd.n78 dvdd 2.9391
R13238 dvdd.n82 dvdd 2.9391
R13239 dvdd.n86 dvdd 2.9391
R13240 dvdd.n90 dvdd 2.9391
R13241 dvdd.n94 dvdd 2.9391
R13242 dvdd.n105 dvdd.n99 2.90005
R13243 dvdd.n141 dvdd.n136 2.63064
R13244 dvdd.n169 dvdd.n126 2.63064
R13245 dvdd.n160 dvdd.n130 2.27995
R13246 dvdd.n171 dvdd.n170 2.10461
R13247 dvdd.n182 dvdd.n179 1.90772
R13248 dvdd.n187 dvdd.n182 1.90772
R13249 dvdd.n181 dvdd.n180 1.90772
R13250 dvdd.n183 dvdd.n181 1.90772
R13251 dvdd.n303 dvdd.n302 1.69386
R13252 dvdd.n159 dvdd.n157 1.2279
R13253 dvdd.n143 dvdd.n137 1.05227
R13254 dvdd.n121 dvdd.n99 0.955857
R13255 dvdd.n106 dvdd.n105 0.705857
R13256 dvdd.n107 dvdd.n106 0.705857
R13257 dvdd.n113 dvdd.n112 0.705857
R13258 dvdd.n112 dvdd.n111 0.705857
R13259 dvdd.n111 dvdd.n98 0.705857
R13260 dvdd.n192 dvdd 0.645031
R13261 dvdd.n114 dvdd.n107 0.529518
R13262 dvdd.n165 dvdd.n164 0.526527
R13263 dvdd.n122 dvdd.n98 0.346482
R13264 dvdd.n115 dvdd.n114 0.3105
R13265 dvdd.n121 dvdd.n120 0.3105
R13266 dvdd.n114 dvdd.n113 0.176839
R13267 dvdd.n265 dvdd 0.121114
R13268 dvdd.n269 dvdd 0.121114
R13269 dvdd.n273 dvdd 0.121114
R13270 dvdd.n277 dvdd 0.121114
R13271 dvdd.n281 dvdd 0.121114
R13272 dvdd.n285 dvdd 0.121114
R13273 dvdd.n289 dvdd 0.121114
R13274 dvdd.n293 dvdd 0.121114
R13275 dvdd.n297 dvdd 0.121114
R13276 dvdd.n301 dvdd 0.121114
R13277 dvdd.n65 dvdd 0.121114
R13278 dvdd.n69 dvdd 0.121114
R13279 dvdd.n73 dvdd 0.121114
R13280 dvdd.n77 dvdd 0.121114
R13281 dvdd.n81 dvdd 0.121114
R13282 dvdd.n85 dvdd 0.121114
R13283 dvdd.n89 dvdd 0.121114
R13284 dvdd.n93 dvdd 0.121114
R13285 dvdd.n97 dvdd 0.121114
R13286 dvdd.n144 dvdd.n143 0.120292
R13287 dvdd.n145 dvdd.n144 0.120292
R13288 dvdd.n145 dvdd.n134 0.120292
R13289 dvdd.n152 dvdd.n134 0.120292
R13290 dvdd.n153 dvdd.n152 0.120292
R13291 dvdd.n154 dvdd.n153 0.120292
R13292 dvdd.n154 dvdd.n131 0.120292
R13293 dvdd.n161 dvdd.n131 0.120292
R13294 dvdd.n162 dvdd.n161 0.120292
R13295 dvdd.n162 dvdd.n127 0.120292
R13296 dvdd.n167 dvdd.n127 0.120292
R13297 dvdd.n168 dvdd.n167 0.120292
R13298 dvdd.n173 dvdd.n172 0.120292
R13299 dvdd.n174 dvdd.n173 0.120292
R13300 dvdd.n174 dvdd.n123 0.120292
R13301 dvdd.n178 dvdd.n123 0.120292
R13302 dvdd.n172 dvdd 0.0603958
R13303 dvdd dvdd.n265 0.0377807
R13304 dvdd.n266 dvdd 0.0377807
R13305 dvdd dvdd.n269 0.0377807
R13306 dvdd.n270 dvdd 0.0377807
R13307 dvdd dvdd.n273 0.0377807
R13308 dvdd.n274 dvdd 0.0377807
R13309 dvdd dvdd.n277 0.0377807
R13310 dvdd.n278 dvdd 0.0377807
R13311 dvdd dvdd.n281 0.0377807
R13312 dvdd.n282 dvdd 0.0377807
R13313 dvdd dvdd.n285 0.0377807
R13314 dvdd.n286 dvdd 0.0377807
R13315 dvdd dvdd.n289 0.0377807
R13316 dvdd.n290 dvdd 0.0377807
R13317 dvdd dvdd.n293 0.0377807
R13318 dvdd.n294 dvdd 0.0377807
R13319 dvdd dvdd.n297 0.0377807
R13320 dvdd.n298 dvdd 0.0377807
R13321 dvdd dvdd.n301 0.0377807
R13322 dvdd dvdd.n65 0.0377807
R13323 dvdd.n66 dvdd 0.0377807
R13324 dvdd dvdd.n69 0.0377807
R13325 dvdd.n70 dvdd 0.0377807
R13326 dvdd dvdd.n73 0.0377807
R13327 dvdd.n74 dvdd 0.0377807
R13328 dvdd dvdd.n77 0.0377807
R13329 dvdd.n78 dvdd 0.0377807
R13330 dvdd dvdd.n81 0.0377807
R13331 dvdd.n82 dvdd 0.0377807
R13332 dvdd dvdd.n85 0.0377807
R13333 dvdd.n86 dvdd 0.0377807
R13334 dvdd dvdd.n89 0.0377807
R13335 dvdd.n90 dvdd 0.0377807
R13336 dvdd dvdd.n93 0.0377807
R13337 dvdd.n94 dvdd 0.0377807
R13338 dvdd dvdd.n97 0.0377807
R13339 dvdd.n168 dvdd 0.0226354
R13340 dvdd dvdd.n178 0.0226354
R13341 ibias_gen_0.vn0.n9 ibias_gen_0.vn0.t19 50.4613
R13342 ibias_gen_0.vn0.n10 ibias_gen_0.vn0.t19 50.4344
R13343 ibias_gen_0.vn0.n1 ibias_gen_0.vn0.n7 49.6079
R13344 ibias_gen_0.vn0.n4 ibias_gen_0.vn0.t3 49.2687
R13345 ibias_gen_0.vn0.n1 ibias_gen_0.vn0.t3 49.1817
R13346 ibias_gen_0.vn0.t1 ibias_gen_0.vn0.n3 48.1029
R13347 ibias_gen_0.vn0.t20 ibias_gen_0.vn0.n9 48.1029
R13348 ibias_gen_0.vn0.n8 ibias_gen_0.vn0.t1 48.1029
R13349 ibias_gen_0.vn0.n10 ibias_gen_0.vn0.t20 48.1029
R13350 ibias_gen_0.vn0.n0 ibias_gen_0.vn0.t13 22.9447
R13351 ibias_gen_0.Mt4 ibias_gen_0.vn0.n2 21.105
R13352 ibias_gen_0.Mt4 ibias_gen_0.vn0.n15 19.6387
R13353 ibias_gen_0.Mt4 ibias_gen_0.vn0.n14 19.6387
R13354 ibias_gen_0.Mt4 ibias_gen_0.vn0.n13 19.6387
R13355 ibias_gen_0.vn0.n0 ibias_gen_0.vn0.n12 19.6387
R13356 ibias_gen_0.Mt4 ibias_gen_0.vn0.n16 19.6387
R13357 ibias_gen_0.vn0.n6 ibias_gen_0.vn0.n5 13.8791
R13358 ibias_gen_0.vn0.n9 ibias_gen_0.vn0.n8 13.7174
R13359 ibias_gen_0.vn0.n0 ibias_gen_0.vn0.n11 12.7887
R13360 ibias_gen_0.vn0.n11 ibias_gen_0.vn0.n3 7.26784
R13361 ibias_gen_0.vn0.n11 ibias_gen_0.vn0.n10 6.45004
R13362 ibias_gen_0.vn0.n7 ibias_gen_0.vn0.t17 5.5395
R13363 ibias_gen_0.vn0.n7 ibias_gen_0.vn0.t18 5.5395
R13364 ibias_gen_0.vn0.n15 ibias_gen_0.vn0.t14 3.3065
R13365 ibias_gen_0.vn0.n15 ibias_gen_0.vn0.t12 3.3065
R13366 ibias_gen_0.vn0.n14 ibias_gen_0.vn0.t11 3.3065
R13367 ibias_gen_0.vn0.n14 ibias_gen_0.vn0.t9 3.3065
R13368 ibias_gen_0.vn0.n13 ibias_gen_0.vn0.t8 3.3065
R13369 ibias_gen_0.vn0.n13 ibias_gen_0.vn0.t7 3.3065
R13370 ibias_gen_0.vn0.n12 ibias_gen_0.vn0.t16 3.3065
R13371 ibias_gen_0.vn0.n12 ibias_gen_0.vn0.t10 3.3065
R13372 ibias_gen_0.vn0.n5 ibias_gen_0.vn0.t2 3.3065
R13373 ibias_gen_0.vn0.n5 ibias_gen_0.vn0.t4 3.3065
R13374 ibias_gen_0.vn0.n2 ibias_gen_0.vn0.t6 3.3065
R13375 ibias_gen_0.vn0.n2 ibias_gen_0.vn0.t0 3.3065
R13376 ibias_gen_0.vn0.n16 ibias_gen_0.vn0.t5 3.3065
R13377 ibias_gen_0.vn0.n16 ibias_gen_0.vn0.t15 3.3065
R13378 ibias_gen_0.Mt4 ibias_gen_0.vn0.n0 2.11628
R13379 ibias_gen_0.vn0.n6 ibias_gen_0.vn0.n4 1.44615
R13380 ibias_gen_0.vn0.n8 ibias_gen_0.vn0.n1 1.30001
R13381 ibias_gen_0.vn0.n4 ibias_gen_0.vn0.n3 1.16626
R13382 ibias_gen_0.vn0.n1 ibias_gen_0.vn0.n6 1.15267
R13383 ibias_gen_0.vp0.n3 ibias_gen_0.vp0.n1 57.7416
R13384 ibias_gen_0.vp0.n8 ibias_gen_0.vp0.t13 50.9767
R13385 ibias_gen_0.vp0.t13 ibias_gen_0.vp0.n6 50.9767
R13386 ibias_gen_0.vp0.n7 ibias_gen_0.vp0.t2 49.8109
R13387 ibias_gen_0.vp0.n0 ibias_gen_0.vp0.t2 49.7239
R13388 ibias_gen_0.vp0.t4 ibias_gen_0.vp0.n9 48.6451
R13389 ibias_gen_0.vp0.t12 ibias_gen_0.vp0.n6 48.6451
R13390 ibias_gen_0.vp0.n10 ibias_gen_0.vp0.t4 48.6451
R13391 ibias_gen_0.vp0.n8 ibias_gen_0.vp0.t12 48.6451
R13392 ibias_gen_0.vp0.n5 ibias_gen_0.vp0.n4 42.4505
R13393 ibias_gen_0.vp0.n3 ibias_gen_0.vp0.n2 42.4505
R13394 ibias_gen_0.vp0.n14 ibias_gen_0.vp0.n13 18.2113
R13395 ibias_gen_0.vp0.n12 ibias_gen_0.vp0.n11 17.2812
R13396 ibias_gen_0.vp0.n10 ibias_gen_0.vp0.n6 13.7361
R13397 ibias_gen_0.vp0.n9 ibias_gen_0.vp0.n8 13.7361
R13398 ibias_gen_0.vp0.n13 ibias_gen_0.vp0.n12 13.3639
R13399 ibias_gen_0.vp0.n4 ibias_gen_0.vp0.t3 5.5395
R13400 ibias_gen_0.vp0.n4 ibias_gen_0.vp0.t5 5.5395
R13401 ibias_gen_0.vp0.n2 ibias_gen_0.vp0.t8 5.5395
R13402 ibias_gen_0.vp0.n2 ibias_gen_0.vp0.t6 5.5395
R13403 ibias_gen_0.vp0.n1 ibias_gen_0.vp0.t11 5.5395
R13404 ibias_gen_0.vp0.n1 ibias_gen_0.vp0.t9 5.5395
R13405 ibias_gen_0.vp0.n13 ibias_gen_0.vp0.n3 3.97054
R13406 ibias_gen_0.vp0.n12 ibias_gen_0.vp0.n0 3.77198
R13407 ibias_gen_0.vp0.n11 ibias_gen_0.vp0.t1 3.3065
R13408 ibias_gen_0.vp0.n11 ibias_gen_0.vp0.t0 3.3065
R13409 ibias_gen_0.vp0.n14 ibias_gen_0.vp0.t10 3.3065
R13410 ibias_gen_0.vp0.t7 ibias_gen_0.vp0.n14 3.3065
R13411 ibias_gen_0.vp0.n7 ibias_gen_0.vp0.n5 1.47061
R13412 ibias_gen_0.vp0.n0 ibias_gen_0.vp0.n10 1.3293
R13413 ibias_gen_0.vp0.n9 ibias_gen_0.vp0.n7 1.16626
R13414 ibias_gen_0.vp0.n0 ibias_gen_0.vp0.n5 1.13637
R13415 ibias_gen_0.vr.n2 ibias_gen_0.vr.n0 21.7373
R13416 ibias_gen_0.vr.n2 ibias_gen_0.vr.n1 20.4114
R13417 ibias_gen_0.vr.t4 ibias_gen_0.vr.n2 17.6029
R13418 ibias_gen_0.vr.n1 ibias_gen_0.vr.t3 3.3065
R13419 ibias_gen_0.vr.n1 ibias_gen_0.vr.t1 3.3065
R13420 ibias_gen_0.vr.n0 ibias_gen_0.vr.t0 3.3065
R13421 ibias_gen_0.vr.n0 ibias_gen_0.vr.t2 3.3065
R13422 ovout.n2 ovout.n0 243.458
R13423 ovout.n2 ovout.n1 205.059
R13424 ovout.n4 ovout.n3 205.059
R13425 ovout.n6 ovout.n5 205.059
R13426 ovout.n8 ovout.n7 205.059
R13427 ovout.n10 ovout.n9 205.059
R13428 ovout.n12 ovout.n11 205.059
R13429 ovout.n14 ovout.n13 205.059
R13430 ovout.n18 ovout.n16 133.534
R13431 ovout.n18 ovout.n17 99.1759
R13432 ovout.n20 ovout.n19 99.1759
R13433 ovout.n22 ovout.n21 99.1759
R13434 ovout.n24 ovout.n23 99.1759
R13435 ovout.n26 ovout.n25 99.1759
R13436 ovout.n28 ovout.n27 99.1759
R13437 ovout ovout.n29 97.4305
R13438 ovout.n4 ovout.n2 38.4005
R13439 ovout.n6 ovout.n4 38.4005
R13440 ovout.n8 ovout.n6 38.4005
R13441 ovout.n10 ovout.n8 38.4005
R13442 ovout.n12 ovout.n10 38.4005
R13443 ovout.n14 ovout.n12 38.4005
R13444 ovout.n20 ovout.n18 34.3584
R13445 ovout.n22 ovout.n20 34.3584
R13446 ovout.n24 ovout.n22 34.3584
R13447 ovout.n26 ovout.n24 34.3584
R13448 ovout.n28 ovout.n26 34.3584
R13449 ovout.n30 ovout.n28 34.3584
R13450 ovout.n13 ovout.t23 26.5955
R13451 ovout.n13 ovout.t30 26.5955
R13452 ovout.n0 ovout.t18 26.5955
R13453 ovout.n0 ovout.t29 26.5955
R13454 ovout.n1 ovout.t21 26.5955
R13455 ovout.n1 ovout.t27 26.5955
R13456 ovout.n3 ovout.t19 26.5955
R13457 ovout.n3 ovout.t25 26.5955
R13458 ovout.n5 ovout.t31 26.5955
R13459 ovout.n5 ovout.t24 26.5955
R13460 ovout.n7 ovout.t17 26.5955
R13461 ovout.n7 ovout.t28 26.5955
R13462 ovout.n9 ovout.t22 26.5955
R13463 ovout.n9 ovout.t16 26.5955
R13464 ovout.n11 ovout.t20 26.5955
R13465 ovout.n11 ovout.t26 26.5955
R13466 ovout.n29 ovout.t15 24.9236
R13467 ovout.n29 ovout.t6 24.9236
R13468 ovout.n16 ovout.t10 24.9236
R13469 ovout.n16 ovout.t5 24.9236
R13470 ovout.n17 ovout.t13 24.9236
R13471 ovout.n17 ovout.t3 24.9236
R13472 ovout.n19 ovout.t11 24.9236
R13473 ovout.n19 ovout.t1 24.9236
R13474 ovout.n21 ovout.t7 24.9236
R13475 ovout.n21 ovout.t0 24.9236
R13476 ovout.n23 ovout.t9 24.9236
R13477 ovout.n23 ovout.t4 24.9236
R13478 ovout.n25 ovout.t14 24.9236
R13479 ovout.n25 ovout.t8 24.9236
R13480 ovout.n27 ovout.t12 24.9236
R13481 ovout.n27 ovout.t2 24.9236
R13482 ovout.n15 ovout.n14 12.6066
R13483 ovout ovout.n30 11.4429
R13484 ovout ovout.n15 5.81868
R13485 ovout.n15 ovout 4.52868
R13486 ovout.n30 ovout 1.74595
R13487 ibias_gen_0.vp.n8 ibias_gen_0.vp.t4 56.5501
R13488 ibias_gen_0.vp.n4 ibias_gen_0.vp.t10 50.9767
R13489 ibias_gen_0.vp.n5 ibias_gen_0.vp.t10 50.9767
R13490 ibias_gen_0.vp.t9 ibias_gen_0.vp.n6 50.9767
R13491 ibias_gen_0.vp.t8 ibias_gen_0.vp.n4 48.6451
R13492 ibias_gen_0.vp.n7 ibias_gen_0.vp.t9 48.6451
R13493 ibias_gen_0.vp.n6 ibias_gen_0.vp.t7 48.6451
R13494 ibias_gen_0.vp.n5 ibias_gen_0.vp.t8 48.6451
R13495 ibias_gen_0.vp.t7 ibias_gen_0.vp.n3 48.6451
R13496 ibias_gen_0.vp.n0 ibias_gen_0.vp.n9 42.5266
R13497 ibias_gen_0.vp.n0 ibias_gen_0.vp.n2 42.4505
R13498 ibias_gen_0.vp.n11 ibias_gen_0.vp.n10 15.1165
R13499 ibias_gen_0.vp.n10 ibias_gen_0.vp.n1 14.8365
R13500 ibias_gen_0.vp.n8 ibias_gen_0.vp.n7 10.5264
R13501 ibias_gen_0.vp.n10 ibias_gen_0.vp.n0 7.57893
R13502 ibias_gen_0.vp.n0 ibias_gen_0.vp.n8 6.28836
R13503 ibias_gen_0.vp.n2 ibias_gen_0.vp.t6 5.5395
R13504 ibias_gen_0.vp.t0 ibias_gen_0.vp.n2 5.5395
R13505 ibias_gen_0.vp.n9 ibias_gen_0.vp.t0 5.5395
R13506 ibias_gen_0.vp.n9 ibias_gen_0.vp.t2 5.5395
R13507 ibias_gen_0.vp.n1 ibias_gen_0.vp.t3 3.3065
R13508 ibias_gen_0.vp.t1 ibias_gen_0.vp.n1 3.3065
R13509 ibias_gen_0.vp.t1 ibias_gen_0.vp.n11 3.3065
R13510 ibias_gen_0.vp.n11 ibias_gen_0.vp.t5 3.3065
R13511 ibias_gen_0.vp.n6 ibias_gen_0.vp.n5 2.33202
R13512 ibias_gen_0.vp.n4 ibias_gen_0.vp.n3 2.33202
R13513 ibias_gen_0.vp.n7 ibias_gen_0.vp.n3 2.33126
R13514 itest itest.n0 45.907
R13515 itest.n0 itest.t0 5.5395
R13516 itest.n0 itest.t1 5.5395
R13517 rstring_mux_0.vtrip10.n2 rstring_mux_0.vtrip10.n0 50.7022
R13518 rstring_mux_0.vtrip10.n3 rstring_mux_0.vtrip10.n2 17.3151
R13519 rstring_mux_0.vtrip10.n2 rstring_mux_0.vtrip10.n1 13.8791
R13520 rstring_mux_0.vtrip10.n3 rstring_mux_0.vtrip10.t5 10.6303
R13521 rstring_mux_0.vtrip10.n0 rstring_mux_0.vtrip10.t4 5.5395
R13522 rstring_mux_0.vtrip10.n0 rstring_mux_0.vtrip10.t3 5.5395
R13523 rstring_mux_0.vtrip10.n1 rstring_mux_0.vtrip10.t0 3.3065
R13524 rstring_mux_0.vtrip10.n1 rstring_mux_0.vtrip10.t1 3.3065
R13525 rstring_mux_0.vtrip10.t2 rstring_mux_0.vtrip10.n3 0.825482
R13526 schmitt_trigger_0.m.n8 schmitt_trigger_0.m.t14 240.764
R13527 schmitt_trigger_0.m.n9 schmitt_trigger_0.m.t16 240.713
R13528 schmitt_trigger_0.m.n10 schmitt_trigger_0.m.t17 240.529
R13529 schmitt_trigger_0.m.n8 schmitt_trigger_0.m.t15 240.349
R13530 schmitt_trigger_0.m.n7 schmitt_trigger_0.m.n5 211.214
R13531 schmitt_trigger_0.m.n3 schmitt_trigger_0.m.n1 207.804
R13532 schmitt_trigger_0.m.n3 schmitt_trigger_0.m.n2 207.585
R13533 schmitt_trigger_0.m.n4 schmitt_trigger_0.m.n0 204.175
R13534 schmitt_trigger_0.m.n7 schmitt_trigger_0.m.n6 204.175
R13535 schmitt_trigger_0.m.n15 schmitt_trigger_0.m.n14 70.9014
R13536 schmitt_trigger_0.m.n13 schmitt_trigger_0.m.n12 70.9014
R13537 schmitt_trigger_0.m.n0 schmitt_trigger_0.m.t5 28.5655
R13538 schmitt_trigger_0.m.n0 schmitt_trigger_0.m.t6 28.5655
R13539 schmitt_trigger_0.m.n6 schmitt_trigger_0.m.t10 28.5655
R13540 schmitt_trigger_0.m.n6 schmitt_trigger_0.m.t9 28.5655
R13541 schmitt_trigger_0.m.n5 schmitt_trigger_0.m.t13 28.5655
R13542 schmitt_trigger_0.m.n5 schmitt_trigger_0.m.t11 28.5655
R13543 schmitt_trigger_0.m.n1 schmitt_trigger_0.m.t3 28.5655
R13544 schmitt_trigger_0.m.n1 schmitt_trigger_0.m.t4 28.5655
R13545 schmitt_trigger_0.m.n2 schmitt_trigger_0.m.t7 28.5655
R13546 schmitt_trigger_0.m.n2 schmitt_trigger_0.m.t0 28.5655
R13547 schmitt_trigger_0.m.n14 schmitt_trigger_0.m.t2 17.4005
R13548 schmitt_trigger_0.m.n14 schmitt_trigger_0.m.t1 17.4005
R13549 schmitt_trigger_0.m.n12 schmitt_trigger_0.m.t12 17.4005
R13550 schmitt_trigger_0.m.n12 schmitt_trigger_0.m.t8 17.4005
R13551 schmitt_trigger_0.m.n10 schmitt_trigger_0.m.n9 12.9318
R13552 schmitt_trigger_0.m.n11 schmitt_trigger_0.m.n7 8.3606
R13553 schmitt_trigger_0.m.n4 schmitt_trigger_0.m.n3 3.62811
R13554 schmitt_trigger_0.m schmitt_trigger_0.m.n4 0.819515
R13555 schmitt_trigger_0.m schmitt_trigger_0.m.n15 0.73133
R13556 schmitt_trigger_0.m.n15 schmitt_trigger_0.m.n13 0.688
R13557 schmitt_trigger_0.m.n11 schmitt_trigger_0.m.n10 0.358635
R13558 schmitt_trigger_0.m.n13 schmitt_trigger_0.m.n11 0.251558
R13559 schmitt_trigger_0.m.n9 schmitt_trigger_0.m.n8 0.0297969
R13560 ibias_gen_0.vp1.n5 ibias_gen_0.vp1.n4 53.0003
R13561 ibias_gen_0.vp1.t15 ibias_gen_0.vp1.n3 49.8109
R13562 ibias_gen_0.vp1.n3 ibias_gen_0.vp1.t13 49.8109
R13563 ibias_gen_0.vp1.t13 ibias_gen_0.vp1.n0 49.7878
R13564 ibias_gen_0.vp1.n0 ibias_gen_0.vp1.t15 49.6053
R13565 ibias_gen_0.vp1 ibias_gen_0.vp1.n6 45.7548
R13566 ibias_gen_0.vp1.n2 ibias_gen_0.vp1.n1 42.4505
R13567 ibias_gen_0.vp1.n9 ibias_gen_0.vp1.n7 18.5825
R13568 ibias_gen_0.vp1.n15 ibias_gen_0.vp1.n14 17.1535
R13569 ibias_gen_0.vp1.n11 ibias_gen_0.vp1.n10 16.3247
R13570 ibias_gen_0.vp1.n9 ibias_gen_0.vp1.n8 16.3247
R13571 ibias_gen_0.vp1.n13 ibias_gen_0.vp1.n12 15.5548
R13572 ibias_gen_0.vp1.n15 ibias_gen_0.vp1.n13 11.684
R13573 ibias_gen_0.vp1.n6 ibias_gen_0.vp1.t0 5.5395
R13574 ibias_gen_0.vp1.n6 ibias_gen_0.vp1.t17 5.5395
R13575 ibias_gen_0.vp1.n4 ibias_gen_0.vp1.t12 5.5395
R13576 ibias_gen_0.vp1.n4 ibias_gen_0.vp1.t2 5.5395
R13577 ibias_gen_0.vp1.n1 ibias_gen_0.vp1.t14 5.5395
R13578 ibias_gen_0.vp1.n1 ibias_gen_0.vp1.t16 5.5395
R13579 ibias_gen_0.vp1.n5 ibias_gen_0.vp1.n0 4.85318
R13580 ibias_gen_0.vp1.n11 ibias_gen_0.vp1.n9 4.51612
R13581 ibias_gen_0.vp1.n12 ibias_gen_0.vp1.t9 3.3065
R13582 ibias_gen_0.vp1.n12 ibias_gen_0.vp1.t4 3.3065
R13583 ibias_gen_0.vp1.n10 ibias_gen_0.vp1.t11 3.3065
R13584 ibias_gen_0.vp1.n10 ibias_gen_0.vp1.t8 3.3065
R13585 ibias_gen_0.vp1.n8 ibias_gen_0.vp1.t7 3.3065
R13586 ibias_gen_0.vp1.n8 ibias_gen_0.vp1.t10 3.3065
R13587 ibias_gen_0.vp1.n7 ibias_gen_0.vp1.t5 3.3065
R13588 ibias_gen_0.vp1.n7 ibias_gen_0.vp1.t6 3.3065
R13589 ibias_gen_0.vp1.n14 ibias_gen_0.vp1.t1 3.3065
R13590 ibias_gen_0.vp1.n14 ibias_gen_0.vp1.t3 3.3065
R13591 ibias_gen_0.vp1.n13 ibias_gen_0.vp1.n11 2.27562
R13592 ibias_gen_0.vp1 ibias_gen_0.vp1.n15 1.87819
R13593 ibias_gen_0.vp1.n2 ibias_gen_0.vp1.n0 1.48628
R13594 ibias_gen_0.vp1.n3 ibias_gen_0.vp1.n2 1.47061
R13595 ibias_gen_0.vp1 ibias_gen_0.vp1.n5 1.36236
R13596 ibias_gen_0.vn1.n0 ibias_gen_0.vn1.n1 47.4959
R13597 ibias_gen_0.vn1.n3 ibias_gen_0.vn1.t14 27.5855
R13598 ibias_gen_0.vn1.n2 ibias_gen_0.vn1.t10 27.5855
R13599 ibias_gen_0.vn1.n6 ibias_gen_0.vn1.t16 27.5855
R13600 ibias_gen_0.vn1.n5 ibias_gen_0.vn1.t12 27.5855
R13601 ibias_gen_0.vn1.n10 ibias_gen_0.vn1.t6 26.004
R13602 ibias_gen_0.vn1.n0 ibias_gen_0.vn1.n13 24.5059
R13603 ibias_gen_0.vn1.n3 ibias_gen_0.vn1.t17 24.3247
R13604 ibias_gen_0.vn1.n2 ibias_gen_0.vn1.t15 24.3247
R13605 ibias_gen_0.vn1.n6 ibias_gen_0.vn1.t13 24.3247
R13606 ibias_gen_0.vn1.n5 ibias_gen_0.vn1.t11 24.3247
R13607 ibias_gen_0.vn1.n9 ibias_gen_0.vn1.t4 24.3247
R13608 ibias_gen_0.vn1.n14 ibias_gen_0.vn1.n0 17.1535
R13609 ibias_gen_0.vn1.n12 ibias_gen_0.vn1.n11 13.8791
R13610 ibias_gen_0.vn1.n0 ibias_gen_0.vn1.n12 12.7397
R13611 ibias_gen_0.vn1.n1 ibias_gen_0.vn1.t9 5.5395
R13612 ibias_gen_0.vn1.n1 ibias_gen_0.vn1.t1 5.5395
R13613 ibias_gen_0.vn1.n4 ibias_gen_0.vn1.n2 4.66645
R13614 ibias_gen_0.vn1.n7 ibias_gen_0.vn1.n5 4.66645
R13615 ibias_gen_0.vn1.n13 ibias_gen_0.vn1.t0 3.3065
R13616 ibias_gen_0.vn1.n13 ibias_gen_0.vn1.t8 3.3065
R13617 ibias_gen_0.vn1.n11 ibias_gen_0.vn1.t5 3.3065
R13618 ibias_gen_0.vn1.n11 ibias_gen_0.vn1.t7 3.3065
R13619 ibias_gen_0.vn1.n14 ibias_gen_0.vn1.t3 3.3065
R13620 ibias_gen_0.vn1.t2 ibias_gen_0.vn1.n14 3.3065
R13621 ibias_gen_0.vn1.n8 ibias_gen_0.vn1.n4 2.41645
R13622 ibias_gen_0.vn1.n8 ibias_gen_0.vn1.n7 2.41645
R13623 ibias_gen_0.vn1.n4 ibias_gen_0.vn1.n3 2.2505
R13624 ibias_gen_0.vn1.n7 ibias_gen_0.vn1.n6 2.2505
R13625 ibias_gen_0.vn1.n9 ibias_gen_0.vn1.n8 2.2505
R13626 ibias_gen_0.vn1.n10 ibias_gen_0.vn1.n9 1.58202
R13627 ibias_gen_0.vn1.n12 ibias_gen_0.vn1.n10 1.37822
R13628 otrip_decoded[11].n0 otrip_decoded[11].t1 186.374
R13629 otrip_decoded[11].n0 otrip_decoded[11].t0 170.308
R13630 otrip_decoded[11] otrip_decoded[11].n1 154.56
R13631 otrip_decoded[11].n2 otrip_decoded[11].n1 153.462
R13632 otrip_decoded[11].n1 otrip_decoded[11].n0 101.513
R13633 otrip_decoded[11].n3 otrip_decoded[11] 11.8005
R13634 otrip_decoded[11].n3 otrip_decoded[11].n2 4.96991
R13635 otrip_decoded[11].n2 otrip_decoded[11] 3.46403
R13636 otrip_decoded[11] otrip_decoded[11].n3 2.71109
R13637 vbg_1v2.n20 vbg_1v2.t22 384.709
R13638 vbg_1v2.t22 vbg_1v2.n19 384.709
R13639 vbg_1v2.t10 vbg_1v2.n30 384.226
R13640 vbg_1v2.n31 vbg_1v2.t10 384.226
R13641 vbg_1v2.n29 vbg_1v2.t25 384.226
R13642 vbg_1v2.t25 vbg_1v2.n16 384.226
R13643 vbg_1v2.n28 vbg_1v2.t1 384.226
R13644 vbg_1v2.t1 vbg_1v2.n27 384.226
R13645 vbg_1v2.t3 vbg_1v2.n17 384.226
R13646 vbg_1v2.n26 vbg_1v2.t3 384.226
R13647 vbg_1v2.t5 vbg_1v2.n24 384.226
R13648 vbg_1v2.n25 vbg_1v2.t5 384.226
R13649 vbg_1v2.n23 vbg_1v2.t12 384.226
R13650 vbg_1v2.t12 vbg_1v2.n18 384.226
R13651 vbg_1v2.n22 vbg_1v2.t15 384.226
R13652 vbg_1v2.t15 vbg_1v2.n21 384.226
R13653 vbg_1v2.t19 vbg_1v2.n19 384.226
R13654 vbg_1v2.n20 vbg_1v2.t19 384.226
R13655 vbg_1v2.t16 vbg_1v2.n15 384.226
R13656 vbg_1v2.n32 vbg_1v2.t16 384.226
R13657 vbg_1v2 vbg_1v2.n14 20.1485
R13658 vbg_1v2.n7 vbg_1v2.t8 16.6244
R13659 vbg_1v2.n0 vbg_1v2.t24 16.4695
R13660 vbg_1v2.n13 vbg_1v2.t21 16.0763
R13661 vbg_1v2.n12 vbg_1v2.t23 16.0763
R13662 vbg_1v2.n11 vbg_1v2.t18 16.0763
R13663 vbg_1v2.n10 vbg_1v2.t20 16.0763
R13664 vbg_1v2.n9 vbg_1v2.t17 16.0763
R13665 vbg_1v2.n8 vbg_1v2.t13 16.0763
R13666 vbg_1v2.n7 vbg_1v2.t14 16.0763
R13667 vbg_1v2.n6 vbg_1v2.t9 15.9214
R13668 vbg_1v2.n5 vbg_1v2.t11 15.9214
R13669 vbg_1v2.n4 vbg_1v2.t6 15.9214
R13670 vbg_1v2.n3 vbg_1v2.t7 15.9214
R13671 vbg_1v2.n2 vbg_1v2.t4 15.9214
R13672 vbg_1v2.n1 vbg_1v2.t0 15.9214
R13673 vbg_1v2.n0 vbg_1v2.t2 15.9214
R13674 vbg_1v2.n14 vbg_1v2.n6 8.60262
R13675 vbg_1v2.n33 vbg_1v2.n15 7.13992
R13676 vbg_1v2.n14 vbg_1v2.n13 5.62204
R13677 vbg_1v2.n33 vbg_1v2.n32 4.5005
R13678 vbg_1v2.n8 vbg_1v2.n7 0.548577
R13679 vbg_1v2.n9 vbg_1v2.n8 0.548577
R13680 vbg_1v2.n10 vbg_1v2.n9 0.548577
R13681 vbg_1v2.n11 vbg_1v2.n10 0.548577
R13682 vbg_1v2.n12 vbg_1v2.n11 0.548577
R13683 vbg_1v2.n13 vbg_1v2.n12 0.548577
R13684 vbg_1v2.n1 vbg_1v2.n0 0.548577
R13685 vbg_1v2.n2 vbg_1v2.n1 0.548577
R13686 vbg_1v2.n3 vbg_1v2.n2 0.548577
R13687 vbg_1v2.n4 vbg_1v2.n3 0.548577
R13688 vbg_1v2.n5 vbg_1v2.n4 0.548577
R13689 vbg_1v2.n6 vbg_1v2.n5 0.548577
R13690 vbg_1v2.n21 vbg_1v2.n20 0.484196
R13691 vbg_1v2.n21 vbg_1v2.n18 0.484196
R13692 vbg_1v2.n25 vbg_1v2.n18 0.484196
R13693 vbg_1v2.n26 vbg_1v2.n25 0.484196
R13694 vbg_1v2.n27 vbg_1v2.n26 0.484196
R13695 vbg_1v2.n27 vbg_1v2.n16 0.484196
R13696 vbg_1v2.n31 vbg_1v2.n16 0.484196
R13697 vbg_1v2.n22 vbg_1v2.n19 0.484196
R13698 vbg_1v2.n23 vbg_1v2.n22 0.484196
R13699 vbg_1v2.n24 vbg_1v2.n23 0.484196
R13700 vbg_1v2.n24 vbg_1v2.n17 0.484196
R13701 vbg_1v2.n28 vbg_1v2.n17 0.484196
R13702 vbg_1v2.n29 vbg_1v2.n28 0.484196
R13703 vbg_1v2.n30 vbg_1v2.n29 0.484196
R13704 vbg_1v2.n32 vbg_1v2.n31 0.459739
R13705 vbg_1v2.n30 vbg_1v2.n15 0.459739
R13706 vbg_1v2 vbg_1v2.n33 0.063
R13707 rstring_mux_0.vtrip11.n2 rstring_mux_0.vtrip11.n0 50.7022
R13708 rstring_mux_0.vtrip11.n2 rstring_mux_0.vtrip11.n1 13.8791
R13709 rstring_mux_0.vtrip11.t0 rstring_mux_0.vtrip11.n3 10.5857
R13710 rstring_mux_0.vtrip11.n3 rstring_mux_0.vtrip11.t1 10.5847
R13711 rstring_mux_0.vtrip11.n3 rstring_mux_0.vtrip11.n2 9.04505
R13712 rstring_mux_0.vtrip11.n0 rstring_mux_0.vtrip11.t2 5.5395
R13713 rstring_mux_0.vtrip11.n0 rstring_mux_0.vtrip11.t3 5.5395
R13714 rstring_mux_0.vtrip11.n1 rstring_mux_0.vtrip11.t5 3.3065
R13715 rstring_mux_0.vtrip11.n1 rstring_mux_0.vtrip11.t4 3.3065
R13716 ibias_gen_0.vstart.n0 ibias_gen_0.vstart.t0 56.685
R13717 ibias_gen_0.vstart.n5 ibias_gen_0.vstart.n3 20.328
R13718 ibias_gen_0.vstart.n0 ibias_gen_0.vstart.n1 20.2356
R13719 ibias_gen_0.vstart.n5 ibias_gen_0.vstart.n4 20.069
R13720 ibias_gen_0.vstart.n0 ibias_gen_0.vstart.n2 20.069
R13721 ibias_gen_0.vstart.n7 ibias_gen_0.vstart.n6 20.069
R13722 ibias_gen_0.vstart.n4 ibias_gen_0.vstart.t10 3.3065
R13723 ibias_gen_0.vstart.n4 ibias_gen_0.vstart.t1 3.3065
R13724 ibias_gen_0.vstart.n3 ibias_gen_0.vstart.t7 3.3065
R13725 ibias_gen_0.vstart.n3 ibias_gen_0.vstart.t4 3.3065
R13726 ibias_gen_0.vstart.n2 ibias_gen_0.vstart.t5 3.3065
R13727 ibias_gen_0.vstart.n2 ibias_gen_0.vstart.t6 3.3065
R13728 ibias_gen_0.vstart.n1 ibias_gen_0.vstart.t2 3.3065
R13729 ibias_gen_0.vstart.n1 ibias_gen_0.vstart.t3 3.3065
R13730 ibias_gen_0.vstart.n7 ibias_gen_0.vstart.t8 3.3065
R13731 ibias_gen_0.vstart.t9 ibias_gen_0.vstart.n7 3.3065
R13732 ibias_gen_0.vstart.n6 ibias_gen_0.vstart.n0 0.280933
R13733 ibias_gen_0.vstart.n6 ibias_gen_0.vstart.n5 0.2449
R13734 rstring_mux_0.vtrip5.n2 rstring_mux_0.vtrip5.n0 50.7022
R13735 rstring_mux_0.vtrip5.n2 rstring_mux_0.vtrip5.n1 13.8791
R13736 rstring_mux_0.vtrip5.t4 rstring_mux_0.vtrip5.n3 10.5857
R13737 rstring_mux_0.vtrip5.n3 rstring_mux_0.vtrip5.t5 10.5847
R13738 rstring_mux_0.vtrip5.n3 rstring_mux_0.vtrip5.n2 8.40849
R13739 rstring_mux_0.vtrip5.n0 rstring_mux_0.vtrip5.t2 5.5395
R13740 rstring_mux_0.vtrip5.n0 rstring_mux_0.vtrip5.t3 5.5395
R13741 rstring_mux_0.vtrip5.n1 rstring_mux_0.vtrip5.t0 3.3065
R13742 rstring_mux_0.vtrip5.n1 rstring_mux_0.vtrip5.t1 3.3065
R13743 rstring_mux_0.vtrip4.n2 rstring_mux_0.vtrip4.n0 50.7022
R13744 rstring_mux_0.vtrip4.n3 rstring_mux_0.vtrip4.n2 17.28
R13745 rstring_mux_0.vtrip4.n2 rstring_mux_0.vtrip4.n1 13.8791
R13746 rstring_mux_0.vtrip4.n3 rstring_mux_0.vtrip4.t3 10.6297
R13747 rstring_mux_0.vtrip4.n0 rstring_mux_0.vtrip4.t4 5.5395
R13748 rstring_mux_0.vtrip4.n0 rstring_mux_0.vtrip4.t5 5.5395
R13749 rstring_mux_0.vtrip4.n1 rstring_mux_0.vtrip4.t2 3.3065
R13750 rstring_mux_0.vtrip4.n1 rstring_mux_0.vtrip4.t1 3.3065
R13751 rstring_mux_0.vtrip4.t0 rstring_mux_0.vtrip4.n3 0.826075
R13752 otrip_decoded[6].n0 otrip_decoded[6].t0 186.374
R13753 otrip_decoded[6].n0 otrip_decoded[6].t1 170.308
R13754 otrip_decoded[6] otrip_decoded[6].n1 154.56
R13755 otrip_decoded[6].n2 otrip_decoded[6].n1 153.462
R13756 otrip_decoded[6].n1 otrip_decoded[6].n0 101.513
R13757 otrip_decoded[6].n3 otrip_decoded[6] 11.8005
R13758 otrip_decoded[6].n3 otrip_decoded[6].n2 4.96991
R13759 otrip_decoded[6].n2 otrip_decoded[6] 3.46403
R13760 otrip_decoded[6] otrip_decoded[6].n3 2.71109
R13761 rstring_mux_0.vtrip13.n2 rstring_mux_0.vtrip13.n0 50.7022
R13762 rstring_mux_0.vtrip13.n2 rstring_mux_0.vtrip13.n1 13.8791
R13763 rstring_mux_0.vtrip13.t2 rstring_mux_0.vtrip13.n3 10.5857
R13764 rstring_mux_0.vtrip13.n3 rstring_mux_0.vtrip13.t3 10.5847
R13765 rstring_mux_0.vtrip13.n3 rstring_mux_0.vtrip13.n2 9.74147
R13766 rstring_mux_0.vtrip13.n0 rstring_mux_0.vtrip13.t1 5.5395
R13767 rstring_mux_0.vtrip13.n0 rstring_mux_0.vtrip13.t0 5.5395
R13768 rstring_mux_0.vtrip13.n1 rstring_mux_0.vtrip13.t5 3.3065
R13769 rstring_mux_0.vtrip13.n1 rstring_mux_0.vtrip13.t4 3.3065
R13770 schmitt_trigger_0.in.n3 schmitt_trigger_0.in.t10 240.778
R13771 schmitt_trigger_0.in.n0 schmitt_trigger_0.in.t4 240.778
R13772 schmitt_trigger_0.in.n3 schmitt_trigger_0.in.t8 240.349
R13773 schmitt_trigger_0.in.n2 schmitt_trigger_0.in.t1 240.349
R13774 schmitt_trigger_0.in.n1 schmitt_trigger_0.in.t11 240.349
R13775 schmitt_trigger_0.in.n0 schmitt_trigger_0.in.t5 240.349
R13776 schmitt_trigger_0.in.n12 schmitt_trigger_0.in.t2 236.423
R13777 schmitt_trigger_0.in.n12 schmitt_trigger_0.in.t3 236.011
R13778 schmitt_trigger_0.in.n10 schmitt_trigger_0.in.n9 28.545
R13779 schmitt_trigger_0.in.n11 schmitt_trigger_0.in.n10 20.6661
R13780 schmitt_trigger_0.in.n10 schmitt_trigger_0.in.t0 5.93425
R13781 schmitt_trigger_0.in schmitt_trigger_0.in.n12 4.93075
R13782 schmitt_trigger_0.in.n11 schmitt_trigger_0.in.n4 4.72087
R13783 schmitt_trigger_0.in.n1 schmitt_trigger_0.in.n0 0.429848
R13784 schmitt_trigger_0.in.n2 schmitt_trigger_0.in.n1 0.429848
R13785 schmitt_trigger_0.in.n4 schmitt_trigger_0.in.n2 0.285826
R13786 schmitt_trigger_0.in schmitt_trigger_0.in.n11 0.216402
R13787 schmitt_trigger_0.in.n4 schmitt_trigger_0.in.n3 0.0956087
R13788 schmitt_trigger_0.in.n5 schmitt_trigger_0.in.t7 0.0791747
R13789 schmitt_trigger_0.in.n6 schmitt_trigger_0.in.n5 0.06865
R13790 schmitt_trigger_0.in.n7 schmitt_trigger_0.in.n6 0.06865
R13791 schmitt_trigger_0.in.n8 schmitt_trigger_0.in.n7 0.06865
R13792 schmitt_trigger_0.in.n9 schmitt_trigger_0.in.n8 0.06865
R13793 schmitt_trigger_0.in.n5 schmitt_trigger_0.in.t14 0.0110247
R13794 schmitt_trigger_0.in.n6 schmitt_trigger_0.in.t12 0.0110247
R13795 schmitt_trigger_0.in.n7 schmitt_trigger_0.in.t6 0.0110247
R13796 schmitt_trigger_0.in.n8 schmitt_trigger_0.in.t13 0.0110247
R13797 schmitt_trigger_0.in.n9 schmitt_trigger_0.in.t9 0.0110247
R13798 otrip_decoded[4].n0 otrip_decoded[4].t0 186.374
R13799 otrip_decoded[4].n0 otrip_decoded[4].t1 170.308
R13800 otrip_decoded[4] otrip_decoded[4].n1 154.56
R13801 otrip_decoded[4].n2 otrip_decoded[4].n1 153.462
R13802 otrip_decoded[4].n1 otrip_decoded[4].n0 101.513
R13803 otrip_decoded[4].n3 otrip_decoded[4] 11.8005
R13804 otrip_decoded[4].n3 otrip_decoded[4].n2 4.96991
R13805 otrip_decoded[4].n2 otrip_decoded[4] 3.46403
R13806 otrip_decoded[4] otrip_decoded[4].n3 2.71109
R13807 otrip_decoded[9].n0 otrip_decoded[9].t1 186.374
R13808 otrip_decoded[9].n0 otrip_decoded[9].t0 170.308
R13809 otrip_decoded[9] otrip_decoded[9].n1 154.56
R13810 otrip_decoded[9].n2 otrip_decoded[9].n1 153.462
R13811 otrip_decoded[9].n1 otrip_decoded[9].n0 101.513
R13812 otrip_decoded[9].n3 otrip_decoded[9] 11.8005
R13813 otrip_decoded[9].n3 otrip_decoded[9].n2 4.96991
R13814 otrip_decoded[9].n2 otrip_decoded[9] 3.46403
R13815 otrip_decoded[9] otrip_decoded[9].n3 2.71109
R13816 rstring_mux_0.vtop.n4 rstring_mux_0.vtop.t17 87.3599
R13817 rstring_mux_0.vtop.n2 rstring_mux_0.vtop.n0 48.5415
R13818 rstring_mux_0.vtop.n13 rstring_mux_0.vtop.n12 48.4284
R13819 rstring_mux_0.vtop.n11 rstring_mux_0.vtop.n10 48.4284
R13820 rstring_mux_0.vtop.n9 rstring_mux_0.vtop.n8 48.4284
R13821 rstring_mux_0.vtop.n7 rstring_mux_0.vtop.n6 48.4284
R13822 rstring_mux_0.vtop.n2 rstring_mux_0.vtop.n1 48.4284
R13823 rstring_mux_0.vtop.n15 rstring_mux_0.vtop.n14 45.0184
R13824 rstring_mux_0.vtop.n4 rstring_mux_0.vtop.n3 45.0184
R13825 rstring_mux_0.vtop rstring_mux_0.vtop.t0 25.3478
R13826 rstring_mux_0.vtop.n14 rstring_mux_0.vtop.t4 5.5395
R13827 rstring_mux_0.vtop.n14 rstring_mux_0.vtop.t11 5.5395
R13828 rstring_mux_0.vtop.n12 rstring_mux_0.vtop.t5 5.5395
R13829 rstring_mux_0.vtop.n12 rstring_mux_0.vtop.t13 5.5395
R13830 rstring_mux_0.vtop.n10 rstring_mux_0.vtop.t7 5.5395
R13831 rstring_mux_0.vtop.n10 rstring_mux_0.vtop.t15 5.5395
R13832 rstring_mux_0.vtop.n8 rstring_mux_0.vtop.t2 5.5395
R13833 rstring_mux_0.vtop.n8 rstring_mux_0.vtop.t9 5.5395
R13834 rstring_mux_0.vtop.n6 rstring_mux_0.vtop.t3 5.5395
R13835 rstring_mux_0.vtop.n6 rstring_mux_0.vtop.t10 5.5395
R13836 rstring_mux_0.vtop.n3 rstring_mux_0.vtop.t14 5.5395
R13837 rstring_mux_0.vtop.n3 rstring_mux_0.vtop.t12 5.5395
R13838 rstring_mux_0.vtop.n1 rstring_mux_0.vtop.t16 5.5395
R13839 rstring_mux_0.vtop.n1 rstring_mux_0.vtop.t6 5.5395
R13840 rstring_mux_0.vtop.n0 rstring_mux_0.vtop.t1 5.5395
R13841 rstring_mux_0.vtop.n0 rstring_mux_0.vtop.t8 5.5395
R13842 rstring_mux_0.vtop.n15 rstring_mux_0.vtop.n13 3.5118
R13843 rstring_mux_0.vtop.n5 rstring_mux_0.vtop.n4 3.4105
R13844 rstring_mux_0.vtop rstring_mux_0.vtop.n15 0.841716
R13845 rstring_mux_0.vtop.n5 rstring_mux_0.vtop.n2 0.113554
R13846 rstring_mux_0.vtop.n7 rstring_mux_0.vtop.n5 0.113554
R13847 rstring_mux_0.vtop.n9 rstring_mux_0.vtop.n7 0.113554
R13848 rstring_mux_0.vtop.n11 rstring_mux_0.vtop.n9 0.113554
R13849 rstring_mux_0.vtop.n13 rstring_mux_0.vtop.n11 0.113554
R13850 rstring_mux_0.vtrip6.n2 rstring_mux_0.vtrip6.n0 50.7022
R13851 rstring_mux_0.vtrip6.n3 rstring_mux_0.vtrip6.n2 16.583
R13852 rstring_mux_0.vtrip6.n2 rstring_mux_0.vtrip6.n1 13.8791
R13853 rstring_mux_0.vtrip6.n3 rstring_mux_0.vtrip6.t3 10.6303
R13854 rstring_mux_0.vtrip6.n0 rstring_mux_0.vtrip6.t5 5.5395
R13855 rstring_mux_0.vtrip6.n0 rstring_mux_0.vtrip6.t4 5.5395
R13856 rstring_mux_0.vtrip6.n1 rstring_mux_0.vtrip6.t1 3.3065
R13857 rstring_mux_0.vtrip6.n1 rstring_mux_0.vtrip6.t0 3.3065
R13858 rstring_mux_0.vtrip6.t2 rstring_mux_0.vtrip6.n3 0.825482
R13859 otrip_decoded[2].n0 otrip_decoded[2].t0 186.374
R13860 otrip_decoded[2].n0 otrip_decoded[2].t1 170.308
R13861 otrip_decoded[2] otrip_decoded[2].n1 154.56
R13862 otrip_decoded[2].n2 otrip_decoded[2].n1 153.462
R13863 otrip_decoded[2].n1 otrip_decoded[2].n0 101.513
R13864 otrip_decoded[2].n3 otrip_decoded[2] 11.8005
R13865 otrip_decoded[2].n3 otrip_decoded[2].n2 4.96991
R13866 otrip_decoded[2].n2 otrip_decoded[2] 3.46403
R13867 otrip_decoded[2] otrip_decoded[2].n3 2.71109
R13868 ibias_gen_0.ve.t3 ibias_gen_0.ve.n0 31281
R13869 ibias_gen_0.ve.n1 ibias_gen_0.ve.t3 146.25
R13870 ibias_gen_0.ve.n5 ibias_gen_0.ve.n4 56.1758
R13871 ibias_gen_0.ve.n4 ibias_gen_0.ve.n3 21.4999
R13872 ibias_gen_0.ve.n4 ibias_gen_0.ve.n2 20.6571
R13873 ibias_gen_0.ve.n5 ibias_gen_0.ve.n1 8.57525
R13874 sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0.Emitter ibias_gen_0.ve.n5 6.71196
R13875 ibias_gen_0.ve.n3 ibias_gen_0.ve.t1 3.3065
R13876 ibias_gen_0.ve.n3 ibias_gen_0.ve.t2 3.3065
R13877 ibias_gen_0.ve.n2 ibias_gen_0.ve.t4 3.3065
R13878 ibias_gen_0.ve.n2 ibias_gen_0.ve.t0 3.3065
R13879 sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0.Emitter ibias_gen_0.ve.n1 1.86379
R13880 rstring_mux_0.vtrip1.n2 rstring_mux_0.vtrip1.n0 50.7022
R13881 rstring_mux_0.vtrip1.n2 rstring_mux_0.vtrip1.n1 13.8791
R13882 rstring_mux_0.vtrip1.t2 rstring_mux_0.vtrip1.n3 10.5857
R13883 rstring_mux_0.vtrip1.n3 rstring_mux_0.vtrip1.t5 10.5847
R13884 rstring_mux_0.vtrip1.n3 rstring_mux_0.vtrip1.n2 9.54084
R13885 rstring_mux_0.vtrip1.n0 rstring_mux_0.vtrip1.t1 5.5395
R13886 rstring_mux_0.vtrip1.n0 rstring_mux_0.vtrip1.t0 5.5395
R13887 rstring_mux_0.vtrip1.n1 rstring_mux_0.vtrip1.t4 3.3065
R13888 rstring_mux_0.vtrip1.n1 rstring_mux_0.vtrip1.t3 3.3065
R13889 rstring_mux_0.vtrip0.n2 rstring_mux_0.vtrip0.n0 50.7022
R13890 rstring_mux_0.vtrip0.n3 rstring_mux_0.vtrip0.n2 18.7108
R13891 rstring_mux_0.vtrip0.n2 rstring_mux_0.vtrip0.n1 13.8791
R13892 rstring_mux_0.vtrip0.n3 rstring_mux_0.vtrip0.t3 10.5739
R13893 rstring_mux_0.vtrip0.n0 rstring_mux_0.vtrip0.t0 5.5395
R13894 rstring_mux_0.vtrip0.n0 rstring_mux_0.vtrip0.t1 5.5395
R13895 rstring_mux_0.vtrip0.n1 rstring_mux_0.vtrip0.t5 3.3065
R13896 rstring_mux_0.vtrip0.n1 rstring_mux_0.vtrip0.t4 3.3065
R13897 rstring_mux_0.vtrip0.t2 rstring_mux_0.vtrip0.n3 0.769662
R13898 rstring_mux_0.vtrip3.n2 rstring_mux_0.vtrip3.n0 50.7022
R13899 rstring_mux_0.vtrip3.n2 rstring_mux_0.vtrip3.n1 13.8791
R13900 rstring_mux_0.vtrip3.t2 rstring_mux_0.vtrip3.n3 10.5857
R13901 rstring_mux_0.vtrip3.n3 rstring_mux_0.vtrip3.t5 10.5847
R13902 rstring_mux_0.vtrip3.n3 rstring_mux_0.vtrip3.n2 8.88656
R13903 rstring_mux_0.vtrip3.n0 rstring_mux_0.vtrip3.t3 5.5395
R13904 rstring_mux_0.vtrip3.n0 rstring_mux_0.vtrip3.t4 5.5395
R13905 rstring_mux_0.vtrip3.n1 rstring_mux_0.vtrip3.t0 3.3065
R13906 rstring_mux_0.vtrip3.n1 rstring_mux_0.vtrip3.t1 3.3065
R13907 rstring_mux_0.vtrip15.n2 rstring_mux_0.vtrip15.n0 50.7022
R13908 rstring_mux_0.vtrip15.n2 rstring_mux_0.vtrip15.n1 13.8791
R13909 rstring_mux_0.vtrip15.t2 rstring_mux_0.vtrip15.n3 10.5857
R13910 rstring_mux_0.vtrip15.n3 rstring_mux_0.vtrip15.t3 10.5847
R13911 rstring_mux_0.vtrip15.n3 rstring_mux_0.vtrip15.n2 10.4513
R13912 rstring_mux_0.vtrip15.n0 rstring_mux_0.vtrip15.t5 5.5395
R13913 rstring_mux_0.vtrip15.n0 rstring_mux_0.vtrip15.t4 5.5395
R13914 rstring_mux_0.vtrip15.n1 rstring_mux_0.vtrip15.t0 3.3065
R13915 rstring_mux_0.vtrip15.n1 rstring_mux_0.vtrip15.t1 3.3065
R13916 rstring_mux_0.vtrip2.n2 rstring_mux_0.vtrip2.n0 50.7022
R13917 rstring_mux_0.vtrip2.n3 rstring_mux_0.vtrip2.n2 17.9781
R13918 rstring_mux_0.vtrip2.n2 rstring_mux_0.vtrip2.n1 13.8791
R13919 rstring_mux_0.vtrip2.n3 rstring_mux_0.vtrip2.t5 10.6303
R13920 rstring_mux_0.vtrip2.n0 rstring_mux_0.vtrip2.t2 5.5395
R13921 rstring_mux_0.vtrip2.n0 rstring_mux_0.vtrip2.t3 5.5395
R13922 rstring_mux_0.vtrip2.n1 rstring_mux_0.vtrip2.t1 3.3065
R13923 rstring_mux_0.vtrip2.n1 rstring_mux_0.vtrip2.t0 3.3065
R13924 rstring_mux_0.vtrip2.t4 rstring_mux_0.vtrip2.n3 0.825482
R13925 rstring_mux_0.vtrip7.n2 rstring_mux_0.vtrip7.n0 50.7022
R13926 rstring_mux_0.vtrip7.n2 rstring_mux_0.vtrip7.n1 13.8791
R13927 rstring_mux_0.vtrip7.t0 rstring_mux_0.vtrip7.n3 10.5857
R13928 rstring_mux_0.vtrip7.n3 rstring_mux_0.vtrip7.t3 10.5847
R13929 rstring_mux_0.vtrip7.n3 rstring_mux_0.vtrip7.n2 7.77564
R13930 rstring_mux_0.vtrip7.n0 rstring_mux_0.vtrip7.t4 5.5395
R13931 rstring_mux_0.vtrip7.n0 rstring_mux_0.vtrip7.t5 5.5395
R13932 rstring_mux_0.vtrip7.n1 rstring_mux_0.vtrip7.t1 3.3065
R13933 rstring_mux_0.vtrip7.n1 rstring_mux_0.vtrip7.t2 3.3065
R13934 rstring_mux_0.vtrip14.n2 rstring_mux_0.vtrip14.n0 50.7022
R13935 rstring_mux_0.vtrip14.n3 rstring_mux_0.vtrip14.n2 18.8397
R13936 rstring_mux_0.vtrip14.n2 rstring_mux_0.vtrip14.n1 13.8791
R13937 rstring_mux_0.vtrip14.n3 rstring_mux_0.vtrip14.t1 10.6297
R13938 rstring_mux_0.vtrip14.n0 rstring_mux_0.vtrip14.t5 5.5395
R13939 rstring_mux_0.vtrip14.n0 rstring_mux_0.vtrip14.t4 5.5395
R13940 rstring_mux_0.vtrip14.n1 rstring_mux_0.vtrip14.t3 3.3065
R13941 rstring_mux_0.vtrip14.n1 rstring_mux_0.vtrip14.t2 3.3065
R13942 rstring_mux_0.vtrip14.t0 rstring_mux_0.vtrip14.n3 0.826075
R13943 otrip_decoded[10].n0 otrip_decoded[10].t1 186.374
R13944 otrip_decoded[10].n0 otrip_decoded[10].t0 170.308
R13945 otrip_decoded[10] otrip_decoded[10].n1 154.56
R13946 otrip_decoded[10].n2 otrip_decoded[10].n1 153.462
R13947 otrip_decoded[10].n1 otrip_decoded[10].n0 101.513
R13948 otrip_decoded[10].n3 otrip_decoded[10] 11.8005
R13949 otrip_decoded[10].n3 otrip_decoded[10].n2 4.96991
R13950 otrip_decoded[10].n2 otrip_decoded[10] 3.46403
R13951 otrip_decoded[10] otrip_decoded[10].n3 2.71109
R13952 isrc_sel.n0 isrc_sel.t1 186.374
R13953 isrc_sel.n0 isrc_sel.t0 170.308
R13954 isrc_sel isrc_sel.n1 154.56
R13955 isrc_sel.n2 isrc_sel.n1 153.462
R13956 isrc_sel.n1 isrc_sel.n0 101.513
R13957 isrc_sel.n3 isrc_sel 11.8005
R13958 isrc_sel.n3 isrc_sel.n2 4.96991
R13959 isrc_sel.n2 isrc_sel 3.46403
R13960 isrc_sel isrc_sel.n3 2.71109
R13961 vl.n5 vl.n4 585
R13962 vl.n4 vl.n3 294.937
R13963 vl.n2 vl.t1 286.887
R13964 vl.t1 vl.n1 286.887
R13965 vl.n0 vl.t0 66.4067
R13966 vl.n4 vl.t2 24.6255
R13967 vl.n1 sky130_fd_sc_hvl__lsbufhv2lv_1_0.X 8.35418
R13968 vl.n5 sky130_fd_sc_hvl__lsbufhv2lv_1_0.X 8.08471
R13969 sky130_fd_sc_hvl__lsbufhv2lv_1_0.X vl.n2 6.19839
R13970 vl.n3 vl.n0 5.58939
R13971 sky130_fd_sc_hvl__lsbufhv2lv_1_0.X vl.n0 4.04261
R13972 vl.n2 sky130_fd_sc_hvl__lsbufhv2lv_1_0.X 3.77313
R13973 sky130_fd_sc_hvl__lsbufhv2lv_1_0.X vl.n5 1.88682
R13974 vl.n1 sky130_fd_sc_hvl__lsbufhv2lv_1_0.X 1.61734
R13975 vl.n3 sky130_fd_sc_hvl__lsbufhv2lv_1_0.X 0.340647
R13976 otrip_decoded[8].n0 otrip_decoded[8].t1 186.374
R13977 otrip_decoded[8].n0 otrip_decoded[8].t0 170.308
R13978 otrip_decoded[8] otrip_decoded[8].n1 154.56
R13979 otrip_decoded[8].n2 otrip_decoded[8].n1 153.462
R13980 otrip_decoded[8].n1 otrip_decoded[8].n0 101.513
R13981 otrip_decoded[8].n3 otrip_decoded[8] 11.8005
R13982 otrip_decoded[8].n3 otrip_decoded[8].n2 4.96991
R13983 otrip_decoded[8].n2 otrip_decoded[8] 3.46403
R13984 otrip_decoded[8] otrip_decoded[8].n3 2.71109
R13985 otrip_decoded[13].n0 otrip_decoded[13].t1 186.374
R13986 otrip_decoded[13].n0 otrip_decoded[13].t0 170.308
R13987 otrip_decoded[13] otrip_decoded[13].n1 154.56
R13988 otrip_decoded[13].n2 otrip_decoded[13].n1 153.462
R13989 otrip_decoded[13].n1 otrip_decoded[13].n0 101.513
R13990 otrip_decoded[13].n3 otrip_decoded[13] 11.8005
R13991 otrip_decoded[13].n3 otrip_decoded[13].n2 4.96991
R13992 otrip_decoded[13].n2 otrip_decoded[13] 3.46403
R13993 otrip_decoded[13] otrip_decoded[13].n3 2.71109
R13994 otrip_decoded[15].n0 otrip_decoded[15].t1 186.374
R13995 otrip_decoded[15].n0 otrip_decoded[15].t0 170.308
R13996 otrip_decoded[15] otrip_decoded[15].n1 154.56
R13997 otrip_decoded[15].n2 otrip_decoded[15].n1 153.462
R13998 otrip_decoded[15].n1 otrip_decoded[15].n0 101.513
R13999 otrip_decoded[15].n3 otrip_decoded[15] 11.8005
R14000 otrip_decoded[15].n3 otrip_decoded[15].n2 4.96991
R14001 otrip_decoded[15].n2 otrip_decoded[15] 3.46403
R14002 otrip_decoded[15] otrip_decoded[15].n3 2.71109
R14003 ena.n0 ena.t1 186.374
R14004 ena.n0 ena.t0 170.308
R14005 ena ena.n1 154.56
R14006 ena.n2 ena.n1 153.462
R14007 ena.n1 ena.n0 101.513
R14008 ena.n3 ena 11.8005
R14009 ena.n3 ena.n2 4.96991
R14010 ena.n2 ena 3.46403
R14011 ena ena.n3 2.71109
R14012 otrip_decoded[12].n0 otrip_decoded[12].t1 186.374
R14013 otrip_decoded[12].n0 otrip_decoded[12].t0 170.308
R14014 otrip_decoded[12] otrip_decoded[12].n1 154.56
R14015 otrip_decoded[12].n2 otrip_decoded[12].n1 153.462
R14016 otrip_decoded[12].n1 otrip_decoded[12].n0 101.513
R14017 otrip_decoded[12].n3 otrip_decoded[12] 11.8005
R14018 otrip_decoded[12].n3 otrip_decoded[12].n2 4.96991
R14019 otrip_decoded[12].n2 otrip_decoded[12] 3.46403
R14020 otrip_decoded[12] otrip_decoded[12].n3 2.71109
R14021 otrip_decoded[7].n0 otrip_decoded[7].t1 186.374
R14022 otrip_decoded[7].n0 otrip_decoded[7].t0 170.308
R14023 otrip_decoded[7] otrip_decoded[7].n1 154.56
R14024 otrip_decoded[7].n2 otrip_decoded[7].n1 153.462
R14025 otrip_decoded[7].n1 otrip_decoded[7].n0 101.513
R14026 otrip_decoded[7].n3 otrip_decoded[7] 11.8005
R14027 otrip_decoded[7].n3 otrip_decoded[7].n2 4.96991
R14028 otrip_decoded[7].n2 otrip_decoded[7] 3.46403
R14029 otrip_decoded[7] otrip_decoded[7].n3 2.71109
R14030 otrip_decoded[14].n0 otrip_decoded[14].t1 186.374
R14031 otrip_decoded[14].n0 otrip_decoded[14].t0 170.308
R14032 otrip_decoded[14] otrip_decoded[14].n1 154.56
R14033 otrip_decoded[14].n2 otrip_decoded[14].n1 153.462
R14034 otrip_decoded[14].n1 otrip_decoded[14].n0 101.513
R14035 otrip_decoded[14].n3 otrip_decoded[14] 11.8005
R14036 otrip_decoded[14].n3 otrip_decoded[14].n2 4.96991
R14037 otrip_decoded[14].n2 otrip_decoded[14] 3.46403
R14038 otrip_decoded[14] otrip_decoded[14].n3 2.71109
R14039 otrip_decoded[5].n0 otrip_decoded[5].t1 186.374
R14040 otrip_decoded[5].n0 otrip_decoded[5].t0 170.308
R14041 otrip_decoded[5] otrip_decoded[5].n1 154.56
R14042 otrip_decoded[5].n2 otrip_decoded[5].n1 153.462
R14043 otrip_decoded[5].n1 otrip_decoded[5].n0 101.513
R14044 otrip_decoded[5].n3 otrip_decoded[5] 11.8005
R14045 otrip_decoded[5].n3 otrip_decoded[5].n2 4.96991
R14046 otrip_decoded[5].n2 otrip_decoded[5] 3.46403
R14047 otrip_decoded[5] otrip_decoded[5].n3 2.71109
R14048 otrip_decoded[3].n0 otrip_decoded[3].t1 186.374
R14049 otrip_decoded[3].n0 otrip_decoded[3].t0 170.308
R14050 otrip_decoded[3] otrip_decoded[3].n1 154.56
R14051 otrip_decoded[3].n2 otrip_decoded[3].n1 153.462
R14052 otrip_decoded[3].n1 otrip_decoded[3].n0 101.513
R14053 otrip_decoded[3].n3 otrip_decoded[3] 11.8005
R14054 otrip_decoded[3].n3 otrip_decoded[3].n2 4.96991
R14055 otrip_decoded[3].n2 otrip_decoded[3] 3.46403
R14056 otrip_decoded[3] otrip_decoded[3].n3 2.71109
R14057 otrip_decoded[1].n0 otrip_decoded[1].t1 186.374
R14058 otrip_decoded[1].n0 otrip_decoded[1].t0 170.308
R14059 otrip_decoded[1] otrip_decoded[1].n1 154.56
R14060 otrip_decoded[1].n2 otrip_decoded[1].n1 153.462
R14061 otrip_decoded[1].n1 otrip_decoded[1].n0 101.513
R14062 otrip_decoded[1].n3 otrip_decoded[1] 11.8005
R14063 otrip_decoded[1].n3 otrip_decoded[1].n2 4.96991
R14064 otrip_decoded[1].n2 otrip_decoded[1] 3.46403
R14065 otrip_decoded[1] otrip_decoded[1].n3 2.71109
C0 a_n6007_n2964# a_n5907_n2876# 0.40546f
C1 a_n16501_n11914# a_n15745_n11914# 0.296258f
C2 a_n26452_n10337# avss 0.476134f
C3 a_n6673_n11914# avss 0.465068f
C4 comparator_0.n0 comparator_0.n1 0.927093f
C5 rstring_mux_0.otrip_decoded_b_avdd[10] avdd 0.903548f
C6 rstring_mux_0.otrip_decoded_avdd[10] avss 1.41004f
C7 a_n25318_n2937# a_n24562_n2937# 0.296258f
C8 a_n3102_n3990# a_n3527_n3946# 0.460766f
C9 a_3748_n1478# rstring_mux_0.otrip_decoded_avdd[11] 0.13699f
C10 a_n5639_n3946# dvdd 0.176016f
C11 a_10874_n1026# avdd 0.17611f
C12 a_4289_n15834# avss 0.466333f
C13 a_n8119_n1230# avdd 0.194982f
C14 ibias_gen_0.ena comparator_0.vn 0.292742f
C15 a_n11965_n11914# avss 0.465068f
C16 rstring_mux_0.otrip_decoded_avdd[14] avdd 1.94965f
C17 a_n8563_n15834# a_n7807_n15834# 0.296258f
C18 a_5423_n11914# a_6179_n11914# 0.296258f
C19 a_n6007_n1230# a_n5907_n1142# 0.40546f
C20 ibias_gen_0.ena itest 0.154848f
C21 rstring_mux_0.otrip_decoded_avdd[11] rstring_mux_0.otrip_decoded_avdd[10] 1.78184f
C22 rstring_mux_0.otrip_decoded_avdd[13] dvdd 0.324463f
C23 a_n4027_n15834# avss 0.466333f
C24 rstring_mux_0.vtop avdd 12.5857f
C25 a_n8119_n2964# otrip_decoded[0] 0.207169f
C26 a_n7751_n3946# avdd 0.143941f
C27 a_n21793_n11914# a_n21037_n11914# 0.296258f
C28 rstring_mux_0.otrip_decoded_b_avdd[5] vin 0.340862f
C29 a_n17257_n11914# avss 0.465505f
C30 a_4553_n1230# otrip_decoded[13] 0.2082f
C31 a_n990_n3990# dvdd 0.104499f
C32 a_n8019_n2876# avdd 0.864385f
C33 comparator_0.vn avdd 0.747837f
C34 a_n8195_9395# avss 0.721623f
C35 a_n12731_9395# a_n11975_9395# 0.296258f
C36 a_2441_n1230# avdd 0.206171f
C37 rstring_mux_0.otrip_decoded_b_avdd[8] avss 0.36282f
C38 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[14] 0.211299f
C39 a_n9319_n15834# avss 0.466333f
C40 avdd itest 0.256348f
C41 dcomp avss 3.70917f
C42 a_n7326_n3990# a_n7751_n3946# 0.460766f
C43 rstring_mux_0.otrip_decoded_avdd[0] rstring_mux_0.otrip_decoded_b_avdd[0] 0.56463f
C44 a_n22549_n11914# avss 0.465068f
C45 a_1122_n2256# avdd 0.607928f
C46 a_n13855_n15834# a_n13099_n15834# 0.296258f
C47 a_4553_n2964# a_4653_n2876# 0.40546f
C48 a_10874_n2222# dvdd 0.468791f
C49 a_n13487_9395# avss 0.460203f
C50 a_n8019_n2876# a_n7326_n3990# 0.264594f
C51 rstring_mux_0.otrip_decoded_avdd[0] vin 0.882514f
C52 a_n22672_n10337# a_n21916_n10337# 0.296258f
C53 ibias_gen_0.ena rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y 0.1256f
C54 avss dvdd 0.110112f
C55 a_n6007_n1230# dvdd 0.385785f
C56 rstring_mux_0.otrip_decoded_avdd[8] avss 1.37856f
C57 a_n14611_n15834# avss 0.466333f
C58 ibias_gen_0.ibias vin 0.45049f
C59 a_9570_n3990# a_9145_n3946# 0.460766f
C60 rstring_mux_0.otrip_decoded_avdd[4] rstring_mux_0.otrip_decoded_b_avdd[4] 0.57199f
C61 a_2541_n2876# avdd 0.863791f
C62 comparator_0.vt avss 21.649801f
C63 a_n27085_n11914# a_n26329_n11914# 0.296258f
C64 a_n3895_n2964# a_n3527_n3946# 0.138963f
C65 a_n27841_n11914# avss 0.468954f
C66 a_n5907_n2876# a_n4700_n3212# 0.28899f
C67 comparator_0.n1 dcomp 1.7035f
C68 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.otrip_decoded_avdd[2] 0.101824f
C69 a_3234_n2256# a_2809_n2212# 0.460766f
C70 rstring_mux_0.otrip_decoded_avdd[12] avdd 1.6421f
C71 a_8777_n1230# a_9145_n2212# 0.138963f
C72 a_n1415_n3946# dvdd 0.176016f
C73 a_8069_n15834# a_8825_n15834# 0.296258f
C74 a_n19903_n15834# avss 0.466333f
C75 rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y avdd 0.839308f
C76 a_4553_n1230# a_4653_n1142# 0.40546f
C77 a_7972_n3212# rstring_mux_0.otrip_decoded_avdd[14] 0.136133f
C78 a_9570_n2256# avdd 0.612302f
C79 a_n8019_n1142# a_n7326_n2256# 0.264594f
C80 a_n10841_1995# avss 0.460203f
C81 rstring_mux_0.otrip_decoded_avdd[9] rstring_mux_0.otrip_decoded_avdd[10] 0.618116f
C82 rstring_mux_0.otrip_decoded_avdd[11] dvdd 0.518093f
C83 a_n6812_n1478# avdd 0.420451f
C84 a_4553_n1230# dvdd 0.379209f
C85 rstring_mux_0.otrip_decoded_avdd[13] rstring_mux_0.otrip_decoded_b_avdd[13] 0.574941f
C86 a_n19147_n15834# a_n18391_n15834# 0.296258f
C87 comparator_0.vnn ibias_gen_0.ibias 1.74645f
C88 ibias_gen_0.ena comparator_0.n0 0.122686f
C89 a_n8185_n11914# a_n7429_n11914# 0.296258f
C90 a_n3102_n3990# dvdd 0.104499f
C91 a_n10085_1995# a_n9329_1995# 0.296258f
C92 rstring_mux_0.otrip_decoded_b_avdd[3] avdd 0.903548f
C93 a_n25195_n15834# avss 0.466333f
C94 a_n5907_n1142# a_n4700_n1478# 0.28899f
C95 a_8777_n2964# ena 0.2082f
C96 a_n23050_n2937# avss 0.474704f
C97 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[12] 0.158489f
C98 a_n3527_n3946# avdd 0.143952f
C99 a_7972_n1478# rstring_mux_0.otrip_decoded_avdd[15] 0.13699f
C100 a_n14999_9395# a_n14243_9395# 0.296258f
C101 a_n6007_n2964# avdd 0.207177f
C102 comparator_0.n0 avdd 0.980591f
C103 a_7691_n11914# avss 0.525451f
C104 a_n990_n2256# avdd 0.607928f
C105 rstring_mux_0.otrip_decoded_b_avdd[10] vin 0.340862f
C106 comparator_0.vt vbg_1v2 18.9966f
C107 a_2777_n15834# a_3533_n15834# 0.296258f
C108 a_3748_n1478# avdd 0.420074f
C109 a_n990_n2256# a_n1415_n2212# 0.460766f
C110 rstring_mux_0.otrip_decoded_avdd[6] avss 1.36421f
C111 a_2441_n1230# a_2809_n2212# 0.138963f
C112 rstring_mux_0.otrip_decoded_b_avdd[13] avss 0.363125f
C113 a_n24439_n15834# a_n23683_n15834# 0.296258f
C114 ibias_gen_0.isrc_sel avss 3.37615f
C115 rstring_mux_0.otrip_decoded_avdd[9] rstring_mux_0.otrip_decoded_b_avdd[8] 0.155269f
C116 a_4653_n2876# a_5860_n3212# 0.28899f
C117 a_n13477_n11914# a_n12721_n11914# 0.296258f
C118 a_n20404_n10337# avss 0.769579f
C119 a_n5639_n2212# dvdd 0.169974f
C120 rstring_mux_0.otrip_decoded_avdd[14] vin 0.880778f
C121 a_n22294_n2937# a_n21538_n2937# 0.296258f
C122 rstring_mux_0.otrip_decoded_avdd[10] avdd 1.70589f
C123 a_4553_n2964# avdd 0.207177f
C124 rstring_mux_0.otrip_decoded_b_avdd[1] avss 0.365652f
C125 a_10337_n15834# avss 0.769026f
C126 rstring_mux_0.otrip_decoded_avdd[9] dvdd 0.336109f
C127 rstring_mux_0.otrip_decoded_avdd[9] rstring_mux_0.otrip_decoded_avdd[8] 1.27145f
C128 a_n5917_n11914# avss 0.465068f
C129 a_n25696_n10337# avss 0.472978f
C130 a_n5539_n15834# a_n4783_n15834# 0.296258f
C131 comparator_0.vn vin 0.723433f
C132 a_2809_n3946# dvdd 0.176016f
C133 a_8447_n11914# a_9203_n11914# 0.296258f
C134 a_4653_n1142# a_5860_n1478# 0.28899f
C135 a_n5214_n3990# dvdd 0.104499f
C136 a_n7751_n2212# avdd 0.142924f
C137 a_n3895_n2964# dvdd 0.380879f
C138 a_n3795_n2876# a_n3102_n3990# 0.264594f
C139 a_5045_n15834# avss 0.466333f
C140 a_n5907_n1142# avdd 0.863296f
C141 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[10] 0.13771f
C142 a_n18769_n11914# a_n18013_n11914# 0.296258f
C143 a_n11209_n11914# avss 0.465068f
C144 a_n5214_n2256# a_n5639_n2212# 0.460766f
C145 rstring_mux_0.otrip_decoded_avdd[12] rstring_mux_0.otrip_decoded_b_avdd[12] 0.572505f
C146 a_n6007_n2964# otrip_decoded[2] 0.2082f
C147 a_n9707_9395# a_n8951_9395# 0.296258f
C148 a_n3102_n2256# avdd 0.607928f
C149 ibias_gen_0.ena dvdd 0.217293f
C150 a_6665_n1230# otrip_decoded[15] 0.2082f
C151 rstring_mux_0.otrip_decoded_b_avdd[8] avdd 0.903548f
C152 comparator_0.vnn comparator_0.vn 0.291123f
C153 rstring_mux_0.otrip_decoded_avdd[4] avss 1.34995f
C154 comparator_0.vpp comparator_0.vm 0.63342f
C155 comparator_0.vt ibias_gen_0.ena 0.275486f
C156 a_697_n3946# avdd 0.143952f
C157 a_n16501_n11914# avss 0.465068f
C158 a_n4700_n3212# avdd 0.421965f
C159 dcomp avdd 6.84083f
C160 a_n3795_n1142# a_n3102_n2256# 0.264594f
C161 a_n10831_n15834# a_n10075_n15834# 0.296258f
C162 a_6665_n2964# dvdd 0.380879f
C163 a_3155_n11914# a_3911_n11914# 0.296258f
C164 a_4653_n1142# avdd 0.863296f
C165 rstring_mux_0.otrip_decoded_avdd[12] vin 0.880779f
C166 a_n8563_n15834# avss 0.466333f
C167 rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y vin 0.340862f
C168 rstring_mux_0.otrip_decoded_avdd[8] avdd 1.64246f
C169 avdd dvdd 38.276302f
C170 a_n24061_n11914# a_n23305_n11914# 0.296258f
C171 a_n21793_n11914# avss 0.465068f
C172 comparator_0.vt avdd 89.9285f
C173 a_n1415_n2212# dvdd 0.169343f
C174 a_n12731_9395# avss 0.460203f
C175 rstring_mux_0.otrip_decoded_avdd[8] rstring_mux_0.otrip_decoded_b_avdd[7] 0.154952f
C176 rstring_mux_0.otrip_decoded_avdd[7] dvdd 0.291878f
C177 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.otrip_decoded_avdd[8] 0.342557f
C178 a_n13855_n15834# avss 0.466333f
C179 rstring_mux_0.otrip_decoded_b_avdd[3] vin 0.340862f
C180 a_5860_n3212# avdd 0.421965f
C181 a_n7326_n3990# dvdd 0.104499f
C182 a_n1783_n2964# a_n1415_n3946# 0.138963f
C183 a_n27085_n11914# avss 0.465096f
C184 a_n16123_n15834# a_n15367_n15834# 0.296258f
C185 rstring_mux_0.otrip_decoded_b_avdd[6] avss 0.36281f
C186 a_n3895_n2964# a_n3795_n2876# 0.40546f
C187 schmitt_trigger_0.in dvdd 2.60999f
C188 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[8] 0.128751f
C189 a_n5161_n11914# a_n4405_n11914# 0.296258f
C190 a_n24940_n10337# a_n24184_n10337# 0.296258f
C191 comparator_0.n0 vin 0.530105f
C192 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.otrip_decoded_b_avdd[3] 0.571961f
C193 a_n19147_n15834# avss 0.466333f
C194 a_7033_n3946# dvdd 0.176016f
C195 comparator_0.vpp avss 1.85492f
C196 ibias_gen_0.ena_b ibias_gen_0.isrc_sel 1.07804f
C197 a_n3527_n2212# avdd 0.142934f
C198 a_n5214_n2256# avdd 0.607928f
C199 a_n10085_1995# avss 0.460203f
C200 a_n3895_n1230# avdd 0.206171f
C201 a_7458_n2256# a_7033_n2212# 0.460766f
C202 rstring_mux_0.otrip_decoded_avdd[2] avss 1.41238f
C203 ibias_gen_0.ena ibias_gen_0.isrc_sel 1.49913f
C204 a_n8119_n1230# otrip_decoded[1] 0.207169f
C205 a_n24439_n15834# avss 0.466333f
C206 a_5801_n15834# a_6557_n15834# 0.296258f
C207 a_n3895_n1230# a_n3795_n1142# 0.40546f
C208 a_n22294_n2937# avss 0.471605f
C209 rstring_mux_0.otrip_decoded_avdd[10] vin 0.88077f
C210 ibias_gen_0.ibias comparator_0.vn 0.590633f
C211 comparator_0.vnn comparator_0.n0 0.42769f
C212 a_4921_n3946# avdd 0.143952f
C213 a_n21415_n15834# a_n20659_n15834# 0.296258f
C214 rstring_mux_0.otrip_decoded_avdd[6] avdd 1.63595f
C215 a_n3795_n2876# avdd 0.863791f
C216 rstring_mux_0.otrip_decoded_b_avdd[13] avdd 0.90363f
C217 a_n10453_n11914# a_n9697_n11914# 0.296258f
C218 ibias_gen_0.vp1 avss 2.07563f
C219 a_8447_n11914# avss 0.525451f
C220 a_429_n2876# a_1122_n3990# 0.264594f
C221 ibias_gen_0.isrc_sel avdd 10.4556f
C222 a_n12353_1995# a_n11597_1995# 0.296258f
C223 a_6665_n1230# avdd 0.206171f
C224 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.otrip_decoded_avdd[6] 1.12965f
C225 rstring_mux_0.otrip_decoded_avdd[5] dvdd 0.426864f
C226 a_4553_n1230# a_4921_n2212# 0.138963f
C227 a_n15479_n3901# ibg_200n 0.401026f
C228 rstring_mux_0.otrip_decoded_b_avdd[1] avdd 0.904297f
C229 a_6665_n2964# a_6765_n2876# 0.40546f
C230 a_2809_n2212# dvdd 0.169343f
C231 comparator_0.vpp vbg_1v2 2.54499f
C232 a_3155_n11914# avss 0.465978f
C233 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[6] 0.105908f
C234 a_n1783_n1230# dvdd 0.385574f
C235 a_6765_n2876# avdd 0.863791f
C236 a_429_n1142# a_1122_n2256# 0.264594f
C237 a_n26707_n15834# a_n25951_n15834# 0.296258f
C238 rstring_mux_0.otrip_decoded_b_avdd[8] vin 0.340862f
C239 a_n7326_n2256# avdd 0.607831f
C240 ibias_gen_0.isrc_sel ibias_gen_0.isrc_sel_b 1.79811f
C241 a_n15745_n11914# a_n14989_n11914# 0.296258f
C242 a_n3795_n2876# a_n2588_n3212# 0.28899f
C243 a_n24940_n10337# avss 0.472978f
C244 a_n5161_n11914# avss 0.475109f
C245 a_n24562_n2937# a_n23806_n2937# 0.296258f
C246 rstring_mux_0.otrip_decoded_b_avdd[11] avss 0.362811f
C247 rstring_mux_0.otrip_decoded_avdd[2] rstring_mux_0.otrip_decoded_b_avdd[2] 0.572197f
C248 comparator_0.ena_b avss 1.7777f
C249 a_6665_n1230# a_6765_n1142# 0.40546f
C250 a_697_n2212# avdd 0.142934f
C251 a_5801_n15834# avss 0.466333f
C252 a_n2588_n1478# avdd 0.420074f
C253 rstring_mux_0.otrip_decoded_avdd[8] vin 0.880783f
C254 a_8777_n1230# dvdd 0.379192f
C255 a_n3895_n2964# otrip_decoded[4] 0.2082f
C256 a_9570_n2256# a_9145_n2212# 0.460766f
C257 a_n10453_n11914# avss 0.465068f
C258 comparator_0.vt vin 18.2264f
C259 a_8777_n1230# isrc_sel 0.2082f
C260 rstring_mux_0.otrip_decoded_avdd[4] avdd 1.53138f
C261 a_n7807_n15834# a_n7051_n15834# 0.296258f
C262 a_6179_n11914# a_6935_n11914# 0.296258f
C263 a_n3795_n1142# a_n2588_n1478# 0.28899f
C264 rstring_mux_0.otrip_decoded_avdd[3] dvdd 0.401793f
C265 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.otrip_decoded_avdd[6] 0.340239f
C266 ibias_gen_0.ibias comparator_0.n0 0.172565f
C267 rstring_mux_0.otrip_decoded_avdd[11] rstring_mux_0.otrip_decoded_b_avdd[11] 0.572316f
C268 a_9145_n3946# avdd 0.143145f
C269 a_n21037_n11914# a_n20281_n11914# 0.296258f
C270 a_n15745_n11914# avss 0.465068f
C271 a_n1783_n2964# avdd 0.207177f
C272 a_7972_n1478# avdd 0.420074f
C273 a_n11975_9395# a_n11219_9395# 0.296258f
C274 a_n7807_n15834# avss 0.466333f
C275 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[4] 0.101976f
C276 ibias_gen_0.ena comparator_0.vpp 0.770707f
C277 comparator_0.vt comparator_0.vnn 4.14025f
C278 a_n21037_n11914# avss 0.465068f
C279 rstring_mux_0.otrip_decoded_avdd[1] avss 1.63066f
C280 a_n2588_n3212# rstring_mux_0.otrip_decoded_avdd[4] 0.1362f
C281 a_n13099_n15834# a_n12343_n15834# 0.296258f
C282 a_6765_n2876# a_7972_n3212# 0.28899f
C283 a_n11975_9395# avss 0.460203f
C284 a_n21916_n10337# a_n21160_n10337# 0.296258f
C285 a_10515_n1026# a_10874_n2222# 0.166612f
C286 rstring_mux_0.otrip_decoded_b_avdd[6] avdd 0.903548f
C287 a_n13099_n15834# avss 0.466333f
C288 a_8777_n2964# avdd 0.207077f
C289 ibias_gen_0.vp1 ibias_gen_0.ena_b 0.142844f
C290 a_329_n2964# a_697_n3946# 0.138963f
C291 a_4653_n2876# a_5346_n3990# 0.264594f
C292 a_n26329_n11914# a_n25573_n11914# 0.296258f
C293 comparator_0.vpp avdd 28.3316f
C294 a_n26329_n11914# avss 0.465068f
C295 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.otrip_decoded_b_avdd[6] 0.155152f
C296 ibias_gen_0.isrc_sel a_n16775_n2223# 0.291728f
C297 rstring_mux_0.otrip_decoded_avdd[6] vin 0.880781f
C298 rstring_mux_0.otrip_decoded_b_avdd[13] vin 0.340862f
C299 ibias_gen_0.ena ibias_gen_0.vp1 0.271659f
C300 rstring_mux_0.otrip_decoded_avdd[2] avdd 1.542f
C301 a_n18391_n15834# avss 0.466333f
C302 a_8825_n15834# a_9581_n15834# 0.296258f
C303 a_n2588_n1478# rstring_mux_0.otrip_decoded_avdd[5] 0.13699f
C304 a_6765_n1142# a_7972_n1478# 0.28899f
C305 a_4921_n2212# avdd 0.142934f
C306 a_n9329_1995# avss 0.460231f
C307 a_329_n2964# dvdd 0.380879f
C308 a_n1683_n1142# avdd 0.863296f
C309 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.otrip_decoded_avdd[4] 1.15427f
C310 a_n18391_n15834# a_n17635_n15834# 0.296258f
C311 a_n6007_n1230# otrip_decoded[3] 0.2082f
C312 sky130_fd_sc_hd__inv_4_0.Y dvdd 1.2747f
C313 a_n27208_n10337# a_n26452_n10337# 0.296258f
C314 rstring_mux_0.otrip_decoded_b_avdd[1] vin 0.342078f
C315 rstring_mux_0.ena_b avss 1.61845f
C316 a_4653_n1142# a_5346_n2256# 0.264594f
C317 a_n7429_n11914# a_n6673_n11914# 0.296258f
C318 a_n23683_n15834# avss 0.466333f
C319 a_n9329_1995# a_n8573_1995# 0.296258f
C320 ibias_gen_0.vp1 avdd 6.78644f
C321 a_n21538_n2937# avss 0.471774f
C322 a_n14621_1995# avss 0.4604f
C323 a_5346_n2256# dvdd 0.104499f
C324 rstring_mux_0.otrip_decoded_b_avdd[4] avss 0.36282f
C325 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[2] 0.10426f
C326 rstring_mux_0.otrip_decoded_avdd[10] rstring_mux_0.otrip_decoded_b_avdd[10] 0.5727f
C327 a_n476_n3212# avdd 0.421965f
C328 rstring_mux_0.otrip_decoded_avdd[0] dvdd 0.197825f
C329 a_9203_n11914# avss 0.525451f
C330 a_8877_n1142# avdd 0.863813f
C331 a_3533_n15834# a_4289_n15834# 0.296258f
C332 ibias_gen_0.ena a_10084_n3212# 0.137017f
C333 a_n26830_n2937# avss 0.787359f
C334 comparator_0.vn comparator_0.n0 1.97882f
C335 comparator_0.vt ibias_gen_0.ibias 0.468817f
C336 ibias_gen_0.ena comparator_0.ena_b 0.707143f
C337 a_n23683_n15834# a_n22927_n15834# 0.296258f
C338 rstring_mux_0.otrip_decoded_avdd[15] avss 1.38048f
C339 a_7458_n3990# dvdd 0.104499f
C340 a_n12721_n11914# a_n11965_n11914# 0.296258f
C341 a_9145_n2212# dvdd 0.169037f
C342 a_3911_n11914# avss 0.484363f
C343 a_n21538_n2937# a_n20782_n2937# 0.296258f
C344 rstring_mux_0.otrip_decoded_avdd[4] vin 0.880782f
C345 a_n14621_1995# a_n13865_1995# 0.296258f
C346 ibias_gen_0.vp1 ibias_gen_0.isrc_sel_b 0.406323f
C347 a_10084_n3212# avdd 0.417292f
C348 a_n8119_n1230# a_n7751_n2212# 0.138963f
C349 rstring_mux_0.otrip_decoded_b_avdd[11] avdd 0.903548f
C350 comparator_0.ena_b avdd 1.00223f
C351 schmitt_trigger_0.in schmitt_trigger_0.m 0.95737f
C352 rstring_mux_0.otrip_decoded_avdd[6] rstring_mux_0.otrip_decoded_b_avdd[5] 0.155092f
C353 a_n1783_n2964# a_n1683_n2876# 0.40546f
C354 a_n4405_n11914# avss 0.482553f
C355 a_n24184_n10337# avss 0.472978f
C356 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.otrip_decoded_avdd[4] 0.503487f
C357 a_n4783_n15834# a_n4027_n15834# 0.296258f
C358 a_5346_n3990# avdd 0.607928f
C359 a_9203_n11914# a_9959_n11914# 0.296258f
C360 ibias_gen_0.isrc_sel a_10084_n1478# 0.155566f
C361 a_n1783_n2964# otrip_decoded[6] 0.2082f
C362 a_7033_n2212# avdd 0.142934f
C363 a_1636_n3212# rstring_mux_0.otrip_decoded_avdd[8] 0.142395f
C364 a_6557_n15834# avss 0.466333f
C365 a_329_n1230# avdd 0.206171f
C366 a_3234_n2256# dvdd 0.104499f
C367 a_n18013_n11914# a_n17257_n11914# 0.296258f
C368 a_n9697_n11914# avss 0.465068f
C369 a_n26830_n2937# a_n26074_n2937# 0.296258f
C370 a_3234_n3990# a_2809_n3946# 0.460766f
C371 ibias_gen_0.ena rstring_mux_0.otrip_decoded_avdd[1] 0.17335f
C372 comparator_0.vm avss 10.3544f
C373 a_n8951_9395# a_n8195_9395# 0.296258f
C374 rstring_mux_0.otrip_decoded_avdd[15] rstring_mux_0.otrip_decoded_b_avdd[14] 0.155139f
C375 a_n1783_n1230# a_n1683_n1142# 0.40546f
C376 rstring_mux_0.otrip_decoded_b_avdd[6] vin 0.340862f
C377 a_10874_n1026# dvdd 0.443515f
C378 a_n8119_n1230# dvdd 0.387414f
C379 comparator_0.vpp vin 1.85152f
C380 a_n14989_n11914# avss 0.465068f
C381 rstring_mux_0.otrip_decoded_b_avdd[9] avss 0.362828f
C382 a_n10075_n15834# a_n9319_n15834# 0.296258f
C383 a_1636_n1478# rstring_mux_0.otrip_decoded_avdd[9] 0.13699f
C384 rstring_mux_0.otrip_decoded_avdd[14] dvdd 0.314216f
C385 a_429_n2876# avdd 0.863791f
C386 rstring_mux_0.otrip_decoded_avdd[13] avss 1.50537f
C387 a_3911_n11914# a_4667_n11914# 0.296258f
C388 rstring_mux_0.otrip_decoded_avdd[1] avdd 1.74762f
C389 rstring_mux_0.otrip_decoded_avdd[2] vin 0.880848f
C390 a_n7051_n15834# avss 0.466333f
C391 a_n23305_n11914# a_n22549_n11914# 0.296258f
C392 a_n7751_n3946# dvdd 0.176029f
C393 a_n20281_n11914# avss 0.465405f
C394 a_10515_n1026# avdd 0.538208f
C395 a_8777_n2964# a_8877_n2876# 0.40546f
C396 a_n11219_9395# avss 0.460203f
C397 rstring_mux_0.vtop a_n27841_n11914# 0.398399f
C398 a_n14243_9395# a_n13487_9395# 0.296258f
C399 a_2441_n1230# dvdd 0.379209f
C400 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.otrip_decoded_avdd[2] 1.42613f
C401 ibias_gen_0.ena rstring_mux_0.ena_b 0.179228f
C402 comparator_0.vt comparator_0.vn 0.201562f
C403 comparator_0.vpp comparator_0.vnn 10.261901f
C404 a_n12343_n15834# avss 0.466333f
C405 a_3234_n3990# avdd 0.607928f
C406 a_n990_n3990# a_n1415_n3946# 0.460766f
C407 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[1] 0.556851f
C408 a_6765_n2876# a_7458_n3990# 0.264594f
C409 a_2441_n2964# a_2809_n3946# 0.138963f
C410 a_n25573_n11914# avss 0.465068f
C411 a_n15367_n15834# a_n14611_n15834# 0.296258f
C412 a_1122_n2256# dvdd 0.104499f
C413 a_n1683_n2876# a_n476_n3212# 0.28899f
C414 a_n24184_n10337# a_n23428_n10337# 0.296258f
C415 a_n4405_n11914# a_n3649_n11914# 0.296258f
C416 a_9570_n3990# avdd 0.60295f
C417 a_n17635_n15834# avss 0.466333f
C418 a_8777_n1230# a_8877_n1142# 0.40546f
C419 rstring_mux_0.ena_b avdd 6.38079f
C420 a_n3895_n1230# otrip_decoded[5] 0.2082f
C421 a_n8119_n2964# avdd 0.194488f
C422 a_n8573_1995# avss 0.4604f
C423 a_1636_n1478# avdd 0.420074f
C424 sky130_fd_sc_hd__inv_4_0.Y ovout 1.46398f
C425 rstring_mux_0.otrip_decoded_b_avdd[4] avdd 0.903548f
C426 ibias_gen_0.ena rstring_mux_0.otrip_decoded_avdd[15] 1.91505f
C427 comparator_0.n1 avss 3.01656f
C428 rstring_mux_0.otrip_decoded_avdd[12] dvdd 0.677007f
C429 a_6557_n15834# a_7313_n15834# 0.296258f
C430 rstring_mux_0.otrip_decoded_avdd[11] avss 1.48249f
C431 a_n22927_n15834# avss 0.466333f
C432 a_n1683_n1142# a_n476_n1478# 0.28899f
C433 rstring_mux_0.otrip_decoded_avdd[14] rstring_mux_0.otrip_decoded_b_avdd[13] 0.155037f
C434 a_n13865_1995# avss 0.460231f
C435 a_n20782_n2937# avss 0.47927f
C436 a_9570_n2256# dvdd 0.103732f
C437 a_n20659_n15834# a_n19903_n15834# 0.296258f
C438 rstring_mux_0.otrip_decoded_b_avdd[11] vin 0.340862f
C439 a_n5214_n3990# a_n5639_n3946# 0.460766f
C440 a_n9697_n11914# a_n8941_n11914# 0.296258f
C441 a_2441_n2964# avdd 0.207177f
C442 a_9959_n11914# avss 0.528805f
C443 a_5860_n3212# rstring_mux_0.otrip_decoded_avdd[12] 0.13761f
C444 rstring_mux_0.otrip_decoded_avdd[15] avdd 1.82f
C445 a_n28219_n15834# avss 0.731654f
C446 a_n11597_1995# a_n10841_1995# 0.296258f
C447 rstring_mux_0.otrip_decoded_b_avdd[14] avss 0.363573f
C448 a_n26074_n2937# avss 0.486052f
C449 comparator_0.n0 dcomp 0.945332f
C450 avss vbg_1v2 6.27979f
C451 rstring_mux_0.otrip_decoded_avdd[9] rstring_mux_0.otrip_decoded_b_avdd[9] 0.572131f
C452 a_1122_n3990# avdd 0.607928f
C453 a_n3527_n3946# dvdd 0.176016f
C454 a_7458_n2256# avdd 0.607928f
C455 a_8877_n2876# a_10084_n3212# 0.28899f
C456 a_4667_n11914# avss 0.525451f
C457 a_n6007_n2964# dvdd 0.380879f
C458 a_n990_n2256# dvdd 0.104499f
C459 rstring_mux_0.otrip_decoded_b_avdd[2] avss 0.363375f
C460 a_n8019_n1142# avdd 0.864468f
C461 a_5346_n2256# a_4921_n2212# 0.460766f
C462 comparator_0.vpp ibias_gen_0.ibias 1.29185f
C463 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[15] 0.377385f
C464 a_5860_n1478# rstring_mux_0.otrip_decoded_avdd[13] 0.13699f
C465 a_n6007_n1230# a_n5639_n2212# 0.138963f
C466 avss ibg_200n 0.598741f
C467 a_n25951_n15834# a_n25195_n15834# 0.296258f
C468 a_n14989_n11914# a_n14233_n11914# 0.296258f
C469 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.otrip_decoded_b_avdd[0] 0.176375f
C470 a_n3649_n11914# avss 0.465525f
C471 a_n23428_n10337# avss 0.472978f
C472 a_329_n2964# otrip_decoded[8] 0.2082f
C473 a_n23806_n2937# a_n23050_n2937# 0.296258f
C474 a_n5639_n3946# avdd 0.145138f
C475 rstring_mux_0.otrip_decoded_avdd[1] vin 0.881159f
C476 a_8877_n1142# a_10084_n1478# 0.28899f
C477 rstring_mux_0.otrip_decoded_avdd[10] dvdd 0.293019f
C478 rstring_mux_0.otrip_decoded_avdd[9] avss 1.39274f
C479 a_n6812_n3212# avdd 0.421965f
C480 comparator_0.vm avdd 0.381919f
C481 a_7313_n15834# avss 0.466333f
C482 a_4553_n2964# dvdd 0.380879f
C483 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.otrip_decoded_b_avdd[4] 0.155007f
C484 a_2541_n1142# avdd 0.863296f
C485 a_n8941_n11914# avss 0.465068f
C486 a_n7051_n15834# a_n6295_n15834# 0.296258f
C487 a_6765_n1142# a_7458_n2256# 0.264594f
C488 a_6935_n11914# a_7691_n11914# 0.296258f
C489 ibias_gen_0.ena_b avss 2.73747f
C490 rstring_mux_0.otrip_decoded_b_avdd[9] avdd 0.903548f
C491 rstring_mux_0.otrip_decoded_avdd[13] avdd 2.25867f
C492 a_n7751_n2212# dvdd 0.169579f
C493 a_1122_n2256# a_697_n2212# 0.460766f
C494 a_n20281_n11914# a_n19525_n11914# 0.296258f
C495 a_n990_n3990# avdd 0.607928f
C496 a_n14233_n11914# avss 0.465264f
C497 a_3748_n3212# avdd 0.421965f
C498 ibias_gen_0.ena avss 14.4989f
C499 a_n5907_n2876# a_n5214_n3990# 0.264594f
C500 a_n11219_9395# a_n10463_9395# 0.296258f
C501 a_n3102_n2256# dvdd 0.104499f
C502 a_n6295_n15834# avss 0.466333f
C503 rstring_mux_0.otrip_decoded_avdd[8] rstring_mux_0.otrip_decoded_b_avdd[8] 0.574058f
C504 a_697_n3946# dvdd 0.176016f
C505 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[13] 0.174324f
C506 a_n19525_n11914# avss 0.467526f
C507 a_10874_n2222# avdd 0.257847f
C508 a_n12343_n15834# a_n11587_n15834# 0.296258f
C509 a_n10463_9395# avss 0.460203f
C510 dcomp dvdd 1.11299f
C511 rstring_mux_0.otrip_decoded_b_avdd[4] vin 0.340862f
C512 avdd avss 2.08641p
C513 a_n21160_n10337# a_n20404_n10337# 0.296258f
C514 a_n6007_n1230# avdd 0.206171f
C515 a_10515_n1026# a_10515_n2156# 0.170258f
C516 comparator_0.vt dcomp 1.45758f
C517 comparator_0.ena_b ibias_gen_0.ibias 0.201288f
C518 a_n11587_n15834# avss 0.466333f
C519 rstring_mux_0.otrip_decoded_b_avdd[7] avss 0.36282f
C520 a_4553_n2964# a_4921_n3946# 0.138963f
C521 a_n25573_n11914# a_n24817_n11914# 0.296258f
C522 a_8877_n2876# a_9570_n3990# 0.264594f
C523 rstring_mux_0.otrip_decoded_avdd[8] dvdd 0.285977f
C524 rstring_mux_0.otrip_decoded_avdd[7] avss 1.37218f
C525 a_n5907_n1142# a_n5214_n2256# 0.264594f
C526 a_n24817_n11914# avss 0.465068f
C527 a_329_n2964# a_429_n2876# 0.40546f
C528 a_n1783_n1230# otrip_decoded[7] 0.2082f
C529 comparator_0.vpp comparator_0.vn 0.326993f
C530 a_n3102_n2256# a_n3527_n2212# 0.460766f
C531 a_n1415_n3946# avdd 0.143952f
C532 a_9581_n15834# a_10337_n15834# 0.296258f
C533 a_n16879_n15834# avss 0.466333f
C534 rstring_mux_0.otrip_decoded_avdd[15] vin 0.880681f
C535 comparator_0.n1 avdd 2.72217f
C536 a_n5907_n2876# avdd 0.863791f
C537 schmitt_trigger_0.in avss 8.07242f
C538 rstring_mux_0.otrip_decoded_avdd[11] avdd 1.88092f
C539 a_4553_n1230# avdd 0.206171f
C540 ibias_gen_0.ena vbg_1v2 0.527591f
C541 rstring_mux_0.otrip_decoded_avdd[4] rstring_mux_0.otrip_decoded_b_avdd[3] 0.155509f
C542 a_n17635_n15834# a_n16879_n15834# 0.296258f
C543 ibias_gen_0.isrc_sel_b avss 2.71097f
C544 a_n26452_n10337# a_n25696_n10337# 0.296258f
C545 a_n6673_n11914# a_n5917_n11914# 0.296258f
C546 a_n3102_n3990# avdd 0.607928f
C547 ibias_gen_0.ena_b ibg_200n 0.467695f
C548 a_n22171_n15834# avss 0.466333f
C549 a_n8573_1995# schmitt_trigger_0.in 0.303942f
C550 a_329_n1230# a_429_n1142# 0.40546f
C551 a_n3527_n2212# dvdd 0.169352f
C552 a_n13109_1995# avss 0.460203f
C553 a_n5214_n2256# dvdd 0.105147f
C554 rstring_mux_0.otrip_decoded_b_avdd[14] avdd 0.904181f
C555 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.otrip_decoded_avdd[0] 3.24722f
C556 a_n3895_n1230# dvdd 0.385808f
C557 ibias_gen_0.ena ibg_200n 0.218863f
C558 avdd vbg_1v2 1.46936f
C559 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[11] 0.14576f
C560 a_4653_n2876# avdd 0.863791f
C561 a_10715_n11914# avss 0.819932f
C562 rstring_mux_0.otrip_decoded_avdd[13] rstring_mux_0.otrip_decoded_b_avdd[12] 0.154961f
C563 a_n27463_n15834# avss 0.466415f
C564 a_4289_n15834# a_5045_n15834# 0.296258f
C565 a_n25318_n2937# avss 0.472952f
C566 rstring_mux_0.otrip_decoded_b_avdd[2] avdd 0.903648f
C567 a_n7326_n2256# a_n7751_n2212# 0.460766f
C568 dcomp ibias_gen_0.isrc_sel 10.963901f
C569 a_n22927_n15834# a_n22171_n15834# 0.296258f
C570 a_n14999_9395# avss 0.721623f
C571 a_4921_n3946# dvdd 0.176016f
C572 rstring_mux_0.otrip_decoded_avdd[6] dvdd 0.258377f
C573 rstring_mux_0.otrip_decoded_avdd[5] avss 1.34873f
C574 a_n5639_n2212# avdd 0.142934f
C575 a_n11965_n11914# a_n11209_n11914# 0.296258f
C576 avdd ibg_200n 0.695438f
C577 a_5423_n11914# avss 0.525451f
C578 a_n4700_n1478# avdd 0.420074f
C579 ibias_gen_0.isrc_sel dvdd 0.174941f
C580 a_n13865_1995# a_n13109_1995# 0.296258f
C581 a_6665_n1230# dvdd 0.379209f
C582 rstring_mux_0.otrip_decoded_b_avdd[9] vin 0.340862f
C583 ibias_gen_0.ena ibias_gen_0.ena_b 1.24167f
C584 rstring_mux_0.otrip_decoded_avdd[13] vin 0.880785f
C585 a_n3895_n1230# a_n3527_n2212# 0.138963f
C586 a_2441_n2964# otrip_decoded[10] 0.2082f
C587 a_n1683_n2876# a_n990_n3990# 0.264594f
C588 rstring_mux_0.otrip_decoded_avdd[9] avdd 1.97541f
C589 a_n22672_n10337# avss 0.472978f
C590 rstring_mux_0.otrip_decoded_b_avdd[12] avss 0.36282f
C591 a_429_n2876# a_1636_n3212# 0.28899f
C592 comparator_0.vpp comparator_0.n0 0.347814f
C593 comparator_0.vnn comparator_0.vm 0.562485f
C594 comparator_0.ena_b comparator_0.vn 1.1214f
C595 a_2809_n3946# avdd 0.143952f
C596 a_9959_n11914# a_10715_n11914# 0.296258f
C597 a_n5214_n3990# avdd 0.607928f
C598 a_n3895_n2964# avdd 0.207177f
C599 a_8069_n15834# avss 0.466333f
C600 a_n28219_n15834# a_n27463_n15834# 0.296258f
C601 ibias_gen_0.ena_b avdd 2.97714f
C602 a_5860_n1478# avdd 0.420074f
C603 rstring_mux_0.otrip_decoded_b_avdd[0] avss 0.399825f
C604 a_n7326_n2256# dvdd 0.104499f
C605 a_n17257_n11914# a_n16501_n11914# 0.296258f
C606 a_n8185_n11914# avss 0.465068f
C607 a_n26074_n2937# a_n25318_n2937# 0.296258f
C608 a_8877_n1142# a_9570_n2256# 0.264594f
C609 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[9] 0.133642f
C610 a_n1683_n1142# a_n990_n2256# 0.264594f
C611 avss vin 18.3765f
C612 ibias_gen_0.ena avdd 13.671599f
C613 a_429_n1142# a_1636_n1478# 0.28899f
C614 a_697_n2212# dvdd 0.169343f
C615 a_2777_n15834# avss 0.466333f
C616 a_n13477_n11914# avss 0.466481f
C617 a_10515_n1026# a_10874_n1026# 0.249533f
C618 a_n9319_n15834# a_n8563_n15834# 0.296258f
C619 a_6665_n2964# avdd 0.207177f
C620 rstring_mux_0.otrip_decoded_avdd[4] dvdd 0.266219f
C621 rstring_mux_0.otrip_decoded_avdd[3] avss 1.341f
C622 a_4667_n11914# a_5423_n11914# 0.296258f
C623 rstring_mux_0.otrip_decoded_avdd[12] rstring_mux_0.otrip_decoded_b_avdd[11] 0.155115f
C624 ibias_gen_0.ena_b ibias_gen_0.isrc_sel_b 3.0701f
C625 a_n5539_n15834# avss 0.466333f
C626 a_n22549_n11914# a_n21793_n11914# 0.296258f
C627 rstring_mux_0.otrip_decoded_avdd[11] vin 0.880778f
C628 a_9145_n3946# dvdd 0.17571f
C629 ibias_gen_0.ena schmitt_trigger_0.in 1.1842f
C630 a_n18769_n11914# avss 0.466224f
C631 comparator_0.vnn avss 2.30923f
C632 a_n1415_n2212# avdd 0.142934f
C633 rstring_mux_0.otrip_decoded_b_avdd[7] avdd 0.903548f
C634 a_n9707_9395# avss 0.460203f
C635 rstring_mux_0.otrip_decoded_avdd[7] avdd 1.82134f
C636 a_n1783_n2964# dvdd 0.380879f
C637 ibias_gen_0.ena ibias_gen_0.isrc_sel_b 1.98919f
C638 a_n3795_n1142# avdd 0.863296f
C639 a_n13487_9395# a_n12731_9395# 0.296258f
C640 a_10874_n2222# a_10515_n2156# 0.249269f
C641 a_n10831_n15834# avss 0.466333f
C642 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.otrip_decoded_b_avdd[7] 0.572384f
C643 a_n7326_n3990# avdd 0.607831f
C644 dvdd ovout 1.54536f
C645 a_329_n1230# otrip_decoded[9] 0.2082f
C646 a_6665_n2964# a_7033_n3946# 0.138963f
C647 a_n24061_n11914# avss 0.465068f
C648 rstring_mux_0.otrip_decoded_b_avdd[14] vin 0.340862f
C649 a_n14611_n15834# a_n13855_n15834# 0.296258f
C650 a_n6812_n3212# rstring_mux_0.otrip_decoded_avdd[0] 0.135767f
C651 schmitt_trigger_0.in avdd 3.97779f
C652 vbg_1v2 vin 5.45404f
C653 a_n23428_n10337# a_n22672_n10337# 0.296258f
C654 ibias_gen_0.ibias comparator_0.vm 0.155234f
C655 a_7033_n3946# avdd 0.143952f
C656 ibias_gen_0.isrc_sel_b avdd 3.34069f
C657 a_n16123_n15834# avss 0.466333f
C658 a_n2588_n3212# avdd 0.421965f
C659 rstring_mux_0.ena_b rstring_mux_0.vtop 2.52783f
C660 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[7] 0.126209f
C661 a_8777_n2964# dvdd 0.38084f
C662 a_n27841_n11914# a_n27085_n11914# 0.296258f
C663 a_n8119_n2964# a_n7751_n3946# 0.138963f
C664 a_n4700_n3212# rstring_mux_0.otrip_decoded_avdd[2] 0.135981f
C665 rstring_mux_0.otrip_decoded_b_avdd[2] vin 0.34139f
C666 a_6765_n1142# avdd 0.863296f
C667 a_n8119_n2964# a_n8019_n2876# 0.40546f
C668 comparator_0.vt comparator_0.vpp 2.58688f
C669 rstring_mux_0.otrip_decoded_b_avdd[5] avss 0.36282f
C670 a_7313_n15834# a_8069_n15834# 0.296258f
C671 a_n21415_n15834# avss 0.466333f
C672 a_n6812_n1478# rstring_mux_0.otrip_decoded_avdd[1] 0.13699f
C673 rstring_mux_0.otrip_decoded_avdd[2] dvdd 0.279505f
C674 a_2541_n2876# a_3234_n3990# 0.264594f
C675 comparator_0.vnn vbg_1v2 2.14732f
C676 a_n12353_1995# avss 0.460203f
C677 a_4921_n2212# dvdd 0.169343f
C678 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.otrip_decoded_b_avdd[2] 0.155546f
C679 rstring_mux_0.otrip_decoded_avdd[15] rstring_mux_0.otrip_decoded_avdd[14] 3.06282f
C680 a_n19903_n15834# a_n19147_n15834# 0.296258f
C681 dcomp ibias_gen_0.vp1 0.654772f
C682 rstring_mux_0.otrip_decoded_avdd[9] vin 0.880777f
C683 a_7972_n3212# avdd 0.421965f
C684 a_n8941_n11914# a_n8185_n11914# 0.296258f
C685 a_n4700_n1478# rstring_mux_0.otrip_decoded_avdd[3] 0.13699f
C686 a_n10841_1995# a_n10085_1995# 0.296258f
C687 a_n26707_n15834# avss 0.466333f
C688 rstring_mux_0.otrip_decoded_avdd[5] avdd 1.83423f
C689 a_n8119_n1230# a_n8019_n1142# 0.40546f
C690 a_n24562_n2937# avss 0.471605f
C691 rstring_mux_0.otrip_decoded_avdd[0] avss 1.64125f
C692 a_2541_n1142# a_3234_n2256# 0.264594f
C693 ibias_gen_0.ibias avss 1.24874f
C694 schmitt_trigger_0.in a_10715_n11914# 0.101853f
C695 a_2809_n2212# avdd 0.142934f
C696 a_6179_n11914# avss 0.525451f
C697 a_n1783_n1230# avdd 0.206171f
C698 a_4553_n2964# otrip_decoded[12] 0.2082f
C699 rstring_mux_0.otrip_decoded_b_avdd[12] avdd 0.903548f
C700 schmitt_trigger_0.m dvdd 2.66806f
C701 ibias_gen_0.ena vin 1.79221f
C702 a_n1783_n1230# a_n1415_n2212# 0.138963f
C703 rstring_mux_0.otrip_decoded_avdd[6] rstring_mux_0.otrip_decoded_b_avdd[6] 0.573474f
C704 a_n25195_n15834# a_n24439_n15834# 0.296258f
C705 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[5] 0.101776f
C706 a_2441_n2964# a_2541_n2876# 0.40546f
C707 a_n14233_n11914# a_n13477_n11914# 0.296258f
C708 a_n21916_n10337# avss 0.472978f
C709 a_n23050_n2937# a_n22294_n2937# 0.296258f
C710 rstring_mux_0.otrip_decoded_b_avdd[0] avdd 0.870606f
C711 a_n16775_n2223# avdd 0.466408f
C712 a_n1683_n2876# avdd 0.863791f
C713 a_8825_n15834# avss 0.466333f
C714 avdd vin 10.6971f
C715 rstring_mux_0.otrip_decoded_avdd[13] rstring_mux_0.otrip_decoded_avdd[14] 1.33995f
C716 a_8777_n1230# avdd 0.206179f
C717 a_n15529_n2223# ibg_200n 0.397003f
C718 a_n8019_n2876# a_n6812_n3212# 0.28899f
C719 a_n7429_n11914# avss 0.465068f
C720 a_n27208_n10337# avss 0.767315f
C721 comparator_0.vn comparator_0.vm 4.6608f
C722 rstring_mux_0.otrip_decoded_avdd[15] rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y 0.572453f
C723 ibias_gen_0.ena comparator_0.vnn 0.738279f
C724 a_n6295_n15834# a_n5539_n15834# 0.296258f
C725 rstring_mux_0.otrip_decoded_b_avdd[7] vin 0.340862f
C726 rstring_mux_0.otrip_decoded_avdd[7] vin 0.880779f
C727 a_7691_n11914# a_8447_n11914# 0.296258f
C728 a_5346_n3990# dvdd 0.104499f
C729 a_2441_n1230# a_2541_n1142# 0.40546f
C730 a_7033_n2212# dvdd 0.169343f
C731 a_3533_n15834# avss 0.466333f
C732 rstring_mux_0.otrip_decoded_avdd[3] avdd 1.95427f
C733 ibias_gen_0.ibias vbg_1v2 1.3306f
C734 rstring_mux_0.otrip_decoded_avdd[2] rstring_mux_0.otrip_decoded_b_avdd[1] 0.155388f
C735 rstring_mux_0.otrip_decoded_b_avdd[10] avss 0.362817f
C736 a_n19525_n11914# a_n18769_n11914# 0.296258f
C737 a_10874_n1026# a_10874_n2222# 0.136815f
C738 a_329_n1230# dvdd 0.379209f
C739 a_n12721_n11914# avss 0.466465f
C740 a_8877_n2876# avdd 0.862949f
C741 ibias_gen_0.vp1 ibias_gen_0.isrc_sel 0.664942f
C742 comparator_0.vnn avdd 28.558f
C743 a_n476_n3212# rstring_mux_0.otrip_decoded_avdd[6] 0.136228f
C744 a_n10463_9395# a_n9707_9395# 0.296258f
C745 a_n8019_n1142# a_n6812_n1478# 0.28899f
C746 ibias_gen_0.ena_b a_n15529_n2223# 0.244191f
C747 a_n4783_n15834# avss 0.466333f
C748 rstring_mux_0.otrip_decoded_avdd[14] avss 1.44633f
C749 a_n18013_n11914# avss 0.466481f
C750 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[3] 0.117254f
C751 a_n11587_n15834# a_n10831_n15834# 0.296258f
C752 rstring_mux_0.otrip_decoded_avdd[11] rstring_mux_0.otrip_decoded_b_avdd[10] 0.155157f
C753 a_n8951_9395# avss 0.460284f
C754 rstring_mux_0.vtop avss 6.96359f
C755 a_n476_n1478# avdd 0.420074f
C756 a_2441_n1230# otrip_decoded[11] 0.2082f
C757 rstring_mux_0.otrip_decoded_avdd[1] dvdd 0.26985f
C758 dcomp a_10515_n1026# 0.207687f
C759 a_n10075_n15834# avss 0.466333f
C760 comparator_0.vn avss 8.805019f
C761 a_n476_n1478# rstring_mux_0.otrip_decoded_avdd[7] 0.13699f
C762 a_n24817_n11914# a_n24061_n11914# 0.296258f
C763 a_8777_n2964# a_9145_n3946# 0.138963f
C764 a_n23305_n11914# avss 0.465068f
C765 a_2541_n2876# a_3748_n3212# 0.28899f
C766 rstring_mux_0.otrip_decoded_avdd[13] rstring_mux_0.otrip_decoded_avdd[12] 2.29107f
C767 a_n14243_9395# avss 0.460284f
C768 a_n15367_n15834# avss 0.466333f
C769 a_5346_n3990# a_4921_n3946# 0.460766f
C770 rstring_mux_0.otrip_decoded_avdd[5] vin 0.880781f
C771 a_3234_n3990# dvdd 0.104499f
C772 a_329_n2964# avdd 0.207177f
C773 rstring_mux_0.otrip_decoded_b_avdd[5] avdd 0.903548f
C774 a_n6007_n2964# a_n5639_n3946# 0.138963f
C775 a_10084_n1478# avdd 0.418567f
C776 ibias_gen_0.ena rstring_mux_0.otrip_decoded_avdd[0] 0.826776f
C777 a_n16879_n15834# a_n16123_n15834# 0.296258f
C778 comparator_0.vm comparator_0.n0 2.59059f
C779 ibias_gen_0.ena ibias_gen_0.ibias 1.6657f
C780 rstring_mux_0.otrip_decoded_avdd[14] rstring_mux_0.otrip_decoded_b_avdd[14] 0.572868f
C781 a_n25696_n10337# a_n24940_n10337# 0.296258f
C782 a_n5917_n11914# a_n5161_n11914# 0.296258f
C783 a_6665_n1230# a_7033_n2212# 0.138963f
C784 a_9570_n3990# dvdd 0.103629f
C785 a_n20659_n15834# avss 0.466333f
C786 a_2541_n1142# a_3748_n1478# 0.28899f
C787 a_5346_n2256# avdd 0.607928f
C788 rstring_mux_0.otrip_decoded_b_avdd[12] vin 0.340862f
C789 a_n8119_n2964# dvdd 0.382499f
C790 a_n11597_1995# avss 0.460203f
C791 rstring_mux_0.otrip_decoded_avdd[12] avss 1.50015f
C792 rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y avss 0.479446f
C793 rstring_mux_0.otrip_decoded_avdd[0] avdd 1.34894f
C794 ibias_gen_0.ibias avdd 2.56431f
C795 a_5045_n15834# a_5801_n15834# 0.296258f
C796 a_n25951_n15834# avss 0.466333f
C797 rstring_mux_0.otrip_decoded_b_avdd[0] vin 0.343304f
C798 a_n23806_n2937# avss 0.474081f
C799 a_7458_n3990# avdd 0.607928f
C800 a_n22171_n15834# a_n21415_n15834# 0.296258f
C801 a_1122_n3990# a_697_n3946# 0.460766f
C802 a_6665_n2964# otrip_decoded[14] 0.2082f
C803 rstring_mux_0.otrip_decoded_b_avdd[3] avss 0.362817f
C804 a_9145_n2212# avdd 0.143323f
C805 a_n11209_n11914# a_n10453_n11914# 0.296258f
C806 a_6935_n11914# avss 0.525451f
C807 a_2441_n2964# dvdd 0.380879f
C808 rstring_mux_0.otrip_decoded_avdd[10] rstring_mux_0.otrip_decoded_b_avdd[9] 0.155018f
C809 a_n13109_1995# a_n12353_1995# 0.296258f
C810 rstring_mux_0.otrip_decoded_avdd[11] rstring_mux_0.otrip_decoded_avdd[12] 1.04751f
C811 a_429_n1142# avdd 0.863296f
C812 rstring_mux_0.otrip_decoded_avdd[15] dvdd 0.289677f
C813 schmitt_trigger_0.in rstring_mux_0.otrip_decoded_avdd[0] 0.260407f
C814 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.otrip_decoded_b_avdd[1] 0.569059f
C815 a_329_n1230# a_697_n2212# 0.138963f
C816 rstring_mux_0.otrip_decoded_avdd[3] vin 0.880782f
C817 comparator_0.n0 avss 3.96407f
C818 a_1122_n3990# dvdd 0.104499f
C819 a_3748_n3212# rstring_mux_0.otrip_decoded_avdd[10] 0.140088f
C820 a_7458_n2256# dvdd 0.104499f
C821 a_n21160_n10337# avss 0.476371f
C822 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.otrip_decoded_b_avdd[5] 0.573322f
C823 a_7458_n3990# a_7033_n3946# 0.460766f
C824 comparator_0.vnn vin 0.772021f
C825 a_1636_n3212# avdd 0.421965f
C826 a_9581_n15834# avss 0.467184f
C827 a_3234_n2256# avdd 0.607928f
C828 a_n27463_n15834# a_n26707_n15834# 0.296258f
C829 ena dvss 0.377679f
C830 otrip_decoded[14] dvss 0.377699f
C831 otrip_decoded[12] dvss 0.377387f
C832 otrip_decoded[10] dvss 0.37758f
C833 otrip_decoded[8] dvss 0.37744f
C834 otrip_decoded[6] dvss 0.378276f
C835 otrip_decoded[4] dvss 0.384187f
C836 otrip_decoded[2] dvss 0.382228f
C837 otrip_decoded[0] dvss 0.403289f
C838 isrc_sel dvss 0.383453f
C839 otrip_decoded[15] dvss 0.375086f
C840 otrip_decoded[13] dvss 0.375086f
C841 otrip_decoded[11] dvss 0.375086f
C842 otrip_decoded[9] dvss 0.375086f
C843 otrip_decoded[7] dvss 0.375086f
C844 otrip_decoded[5] dvss 0.375086f
C845 otrip_decoded[3] dvss 0.374839f
C846 otrip_decoded[1] dvss 0.397873f
C847 ovout dvss 1.33781f
C848 ibg_200n dvss 0.16009f
C849 itest dvss 0.300378f
C850 vin dvss 26.864939f
C851 vbg_1v2 dvss 19.61792f
C852 dvdd dvss 0.181259p
C853 avss dvss 0.165779p
C854 avdd dvss 2.722651p
C855 a_10715_n11914# dvss 0.518783f
C856 a_10337_n15834# dvss 0.542688f
C857 a_9959_n11914# dvss 0.597483f
C858 a_9581_n15834# dvss 0.654446f
C859 a_9203_n11914# dvss 0.659772f
C860 a_8825_n15834# dvss 0.659723f
C861 a_8447_n11914# dvss 0.659772f
C862 a_8069_n15834# dvss 0.659723f
C863 a_7691_n11914# dvss 0.659772f
C864 a_7313_n15834# dvss 0.659723f
C865 a_6935_n11914# dvss 0.659772f
C866 a_6557_n15834# dvss 0.659723f
C867 a_6179_n11914# dvss 0.659772f
C868 a_5801_n15834# dvss 0.659723f
C869 a_5423_n11914# dvss 0.659772f
C870 a_5045_n15834# dvss 0.659723f
C871 a_4667_n11914# dvss 0.659772f
C872 a_4289_n15834# dvss 0.659723f
C873 a_3911_n11914# dvss 0.646333f
C874 a_3533_n15834# dvss 0.644774f
C875 a_3155_n11914# dvss 0.648495f
C876 a_2777_n15834# dvss 0.659723f
C877 a_n3649_n11914# dvss 0.650608f
C878 a_n4027_n15834# dvss 0.659723f
C879 a_n4405_n11914# dvss 0.65628f
C880 a_n4783_n15834# dvss 0.659723f
C881 a_n5161_n11914# dvss 0.659772f
C882 a_n5539_n15834# dvss 0.659723f
C883 a_n5917_n11914# dvss 0.659772f
C884 a_n6295_n15834# dvss 0.659723f
C885 a_n6673_n11914# dvss 0.659772f
C886 a_n7051_n15834# dvss 0.659723f
C887 a_n7429_n11914# dvss 0.659772f
C888 a_n7807_n15834# dvss 0.659723f
C889 a_n8185_n11914# dvss 0.659772f
C890 a_n8563_n15834# dvss 0.659723f
C891 a_n8941_n11914# dvss 0.646141f
C892 a_n9319_n15834# dvss 0.644772f
C893 a_n9697_n11914# dvss 0.658346f
C894 a_n10075_n15834# dvss 0.659723f
C895 a_n10453_n11914# dvss 0.659772f
C896 a_n10831_n15834# dvss 0.659723f
C897 a_n11209_n11914# dvss 0.659772f
C898 a_n11587_n15834# dvss 0.659723f
C899 a_n11965_n11914# dvss 0.659772f
C900 a_n12343_n15834# dvss 0.659723f
C901 a_n12721_n11914# dvss 0.659772f
C902 a_n13099_n15834# dvss 0.659723f
C903 a_n13477_n11914# dvss 0.659772f
C904 a_n13855_n15834# dvss 0.659723f
C905 a_n14233_n11914# dvss 0.659772f
C906 a_n14611_n15834# dvss 0.659723f
C907 a_n14989_n11914# dvss 0.659772f
C908 a_n15367_n15834# dvss 0.645311f
C909 a_n15745_n11914# dvss 0.644801f
C910 a_n16123_n15834# dvss 0.659143f
C911 a_n16501_n11914# dvss 0.659772f
C912 a_n16879_n15834# dvss 0.659723f
C913 a_n17257_n11914# dvss 0.659772f
C914 a_n17635_n15834# dvss 0.659723f
C915 a_n18013_n11914# dvss 0.659772f
C916 a_n18391_n15834# dvss 0.659723f
C917 a_n18769_n11914# dvss 0.659772f
C918 a_n19147_n15834# dvss 0.659723f
C919 a_n19525_n11914# dvss 0.659772f
C920 a_n19903_n15834# dvss 0.659723f
C921 a_n20281_n11914# dvss 0.659772f
C922 a_n20659_n15834# dvss 0.659723f
C923 a_n21037_n11914# dvss 0.659772f
C924 a_n21415_n15834# dvss 0.659723f
C925 a_n21793_n11914# dvss 0.6448f
C926 a_n22171_n15834# dvss 0.644769f
C927 a_n22549_n11914# dvss 0.659772f
C928 a_n22927_n15834# dvss 0.659723f
C929 a_n23305_n11914# dvss 0.659772f
C930 a_n23683_n15834# dvss 0.659723f
C931 a_n24061_n11914# dvss 0.659772f
C932 a_n24439_n15834# dvss 0.659723f
C933 a_n24817_n11914# dvss 0.659772f
C934 a_n25195_n15834# dvss 0.659723f
C935 a_n25573_n11914# dvss 0.659772f
C936 a_n25951_n15834# dvss 0.659723f
C937 a_n26329_n11914# dvss 0.659772f
C938 a_n26707_n15834# dvss 0.659723f
C939 a_n27085_n11914# dvss 0.659772f
C940 a_n27463_n15834# dvss 0.659723f
C941 a_n27841_n11914# dvss 0.659386f
C942 a_n28219_n15834# dvss 0.614933f
C943 rstring_mux_0.vtop dvss 31.8044f
C944 rstring_mux_0.ena_b dvss 2.13314f
C945 rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].Y dvss 0.214336f
C946 rstring_mux_0.otrip_decoded_b_avdd[14] dvss 0.191802f
C947 rstring_mux_0.otrip_decoded_b_avdd[13] dvss 0.191802f
C948 rstring_mux_0.otrip_decoded_b_avdd[12] dvss 0.191802f
C949 rstring_mux_0.otrip_decoded_b_avdd[11] dvss 0.191802f
C950 rstring_mux_0.otrip_decoded_b_avdd[10] dvss 0.191802f
C951 rstring_mux_0.otrip_decoded_b_avdd[9] dvss 0.191801f
C952 rstring_mux_0.otrip_decoded_b_avdd[8] dvss 0.191802f
C953 rstring_mux_0.otrip_decoded_b_avdd[7] dvss 0.191802f
C954 rstring_mux_0.otrip_decoded_b_avdd[6] dvss 0.191802f
C955 rstring_mux_0.otrip_decoded_b_avdd[5] dvss 0.191802f
C956 rstring_mux_0.otrip_decoded_b_avdd[4] dvss 0.191802f
C957 rstring_mux_0.otrip_decoded_b_avdd[3] dvss 0.181122f
C958 rstring_mux_0.otrip_decoded_b_avdd[2] dvss 0.191802f
C959 rstring_mux_0.otrip_decoded_b_avdd[1] dvss 0.191802f
C960 rstring_mux_0.otrip_decoded_b_avdd[0] dvss 0.195093f
C961 a_9145_n3946# dvss 1.71049f
C962 a_7033_n3946# dvss 1.70837f
C963 a_4921_n3946# dvss 1.70837f
C964 a_2809_n3946# dvss 1.70837f
C965 a_697_n3946# dvss 1.70837f
C966 a_n1415_n3946# dvss 1.70837f
C967 a_n3527_n3946# dvss 1.70837f
C968 a_n5639_n3946# dvss 1.70837f
C969 a_n7751_n3946# dvss 1.70982f
C970 a_9570_n3990# dvss 0.891511f
C971 a_7458_n3990# dvss 0.867563f
C972 a_5346_n3990# dvss 0.867563f
C973 rstring_mux_0.otrip_decoded_avdd[14] dvss 1.58527f
C974 a_3234_n3990# dvss 0.867563f
C975 rstring_mux_0.otrip_decoded_avdd[12] dvss 1.58861f
C976 a_1122_n3990# dvss 0.867563f
C977 rstring_mux_0.otrip_decoded_avdd[10] dvss 1.88344f
C978 a_n990_n3990# dvss 0.867563f
C979 rstring_mux_0.otrip_decoded_avdd[8] dvss 1.65793f
C980 a_n3102_n3990# dvss 0.867563f
C981 rstring_mux_0.otrip_decoded_avdd[6] dvss 1.33074f
C982 a_n5214_n3990# dvss 0.867563f
C983 rstring_mux_0.otrip_decoded_avdd[4] dvss 1.07495f
C984 a_n7326_n3990# dvss 0.867659f
C985 rstring_mux_0.otrip_decoded_avdd[2] dvss 1.63868f
C986 rstring_mux_0.otrip_decoded_avdd[0] dvss 1.08019f
C987 a_10084_n3212# dvss 0.508017f
C988 a_8877_n2876# dvss 1.52653f
C989 a_8777_n2964# dvss 1.97982f
C990 a_7972_n3212# dvss 0.503164f
C991 a_6765_n2876# dvss 1.52226f
C992 a_6665_n2964# dvss 1.97975f
C993 a_5860_n3212# dvss 0.503164f
C994 a_4653_n2876# dvss 1.52226f
C995 a_4553_n2964# dvss 1.97975f
C996 a_3748_n3212# dvss 0.503164f
C997 a_2541_n2876# dvss 1.52226f
C998 a_2441_n2964# dvss 1.97975f
C999 a_1636_n3212# dvss 0.503164f
C1000 a_429_n2876# dvss 1.52226f
C1001 a_329_n2964# dvss 1.97975f
C1002 a_n476_n3212# dvss 0.503164f
C1003 a_n1683_n2876# dvss 1.52226f
C1004 a_n1783_n2964# dvss 1.97975f
C1005 a_n2588_n3212# dvss 0.503164f
C1006 a_n3795_n2876# dvss 1.52226f
C1007 a_n3895_n2964# dvss 1.97975f
C1008 a_n4700_n3212# dvss 0.503164f
C1009 a_n5907_n2876# dvss 1.52226f
C1010 a_n6007_n2964# dvss 1.97975f
C1011 a_n6812_n3212# dvss 0.503164f
C1012 a_n8019_n2876# dvss 1.53095f
C1013 a_n8119_n2964# dvss 2.03637f
C1014 a_9145_n2212# dvss 1.69093f
C1015 a_7033_n2212# dvss 1.69148f
C1016 a_10515_n2156# dvss 0.902568f
C1017 a_4921_n2212# dvss 1.69148f
C1018 a_2809_n2212# dvss 1.69148f
C1019 a_697_n2212# dvss 1.69148f
C1020 a_n1415_n2212# dvss 1.69148f
C1021 a_n3527_n2212# dvss 1.69147f
C1022 a_n5639_n2212# dvss 1.69215f
C1023 a_n7751_n2212# dvss 1.69294f
C1024 a_10874_n2222# dvss 1.01173f
C1025 a_9570_n2256# dvss 0.84998f
C1026 a_7458_n2256# dvss 0.867563f
C1027 a_10874_n1026# dvss 0.862185f
C1028 a_10515_n1026# dvss 1.27944f
C1029 a_5346_n2256# dvss 0.867563f
C1030 rstring_mux_0.otrip_decoded_avdd[15] dvss 2.19992f
C1031 a_3234_n2256# dvss 0.867563f
C1032 rstring_mux_0.otrip_decoded_avdd[13] dvss 1.9668f
C1033 a_1122_n2256# dvss 0.867563f
C1034 rstring_mux_0.otrip_decoded_avdd[11] dvss 2.03915f
C1035 a_n990_n2256# dvss 0.867563f
C1036 rstring_mux_0.otrip_decoded_avdd[9] dvss 2.141f
C1037 a_n3102_n2256# dvss 0.867563f
C1038 rstring_mux_0.otrip_decoded_avdd[7] dvss 1.89764f
C1039 a_n5214_n2256# dvss 0.868119f
C1040 rstring_mux_0.otrip_decoded_avdd[5] dvss 2.0224f
C1041 a_n7326_n2256# dvss 0.867659f
C1042 rstring_mux_0.otrip_decoded_avdd[3] dvss 2.12353f
C1043 rstring_mux_0.otrip_decoded_avdd[1] dvss 1.80627f
C1044 a_10084_n1478# dvss 0.490437f
C1045 a_8877_n1142# dvss 1.52856f
C1046 a_8777_n1230# dvss 1.97228f
C1047 a_7972_n1478# dvss 0.501383f
C1048 a_6765_n1142# dvss 1.52953f
C1049 a_6665_n1230# dvss 1.97335f
C1050 a_5860_n1478# dvss 0.501383f
C1051 a_4653_n1142# dvss 1.52953f
C1052 a_4553_n1230# dvss 1.97335f
C1053 a_3748_n1478# dvss 0.501383f
C1054 a_2541_n1142# dvss 1.52953f
C1055 a_2441_n1230# dvss 1.97335f
C1056 a_1636_n1478# dvss 0.501383f
C1057 a_429_n1142# dvss 1.52953f
C1058 a_329_n1230# dvss 1.97335f
C1059 a_n476_n1478# dvss 0.501383f
C1060 a_n1683_n1142# dvss 1.52953f
C1061 a_n1783_n1230# dvss 1.96748f
C1062 a_n2588_n1478# dvss 0.500131f
C1063 a_n3795_n1142# dvss 1.52677f
C1064 a_n3895_n1230# dvss 1.96719f
C1065 a_n4700_n1478# dvss 0.509537f
C1066 a_n5907_n1142# dvss 1.53795f
C1067 a_n6007_n1230# dvss 1.97335f
C1068 a_n6812_n1478# dvss 0.501043f
C1069 a_n8019_n1142# dvss 1.53771f
C1070 a_n8119_n1230# dvss 2.02842f
C1071 sky130_fd_sc_hd__inv_4_0.Y dvss 2.06269f
C1072 schmitt_trigger_0.m dvss 2.476603f
C1073 a_n20404_n10337# dvss 0.639031f
C1074 a_n20782_n2937# dvss 0.502711f
C1075 a_n21160_n10337# dvss 0.639742f
C1076 a_n21538_n2937# dvss 0.502711f
C1077 a_n21916_n10337# dvss 0.646835f
C1078 a_n22294_n2937# dvss 0.502711f
C1079 a_n22672_n10337# dvss 0.639742f
C1080 a_n23050_n2937# dvss 0.502711f
C1081 a_n23428_n10337# dvss 0.639742f
C1082 a_n23806_n2937# dvss 0.502711f
C1083 a_n24184_n10337# dvss 0.639742f
C1084 a_n24562_n2937# dvss 0.502711f
C1085 a_n24940_n10337# dvss 0.639742f
C1086 a_n25318_n2937# dvss 0.502711f
C1087 a_n25696_n10337# dvss 0.639742f
C1088 a_n26074_n2937# dvss 0.502711f
C1089 a_n26452_n10337# dvss 0.639742f
C1090 a_n26830_n2937# dvss 0.502711f
C1091 a_n27208_n10337# dvss 0.638935f
C1092 ibias_gen_0.isrc_sel_b dvss 1.34226f
C1093 ibias_gen_0.isrc_sel dvss 5.29867f
C1094 ibias_gen_0.ena_b dvss 1.24326f
C1095 ibias_gen_0.vp1 dvss 4.856841f
C1096 schmitt_trigger_0.in dvss 0.405956p
C1097 a_n8195_9395# dvss 0.502711f
C1098 a_n8573_1995# dvss 0.502711f
C1099 a_n8951_9395# dvss 0.502711f
C1100 a_n9329_1995# dvss 0.502711f
C1101 a_n9707_9395# dvss 0.502711f
C1102 a_n10085_1995# dvss 0.502711f
C1103 a_n10463_9395# dvss 0.502711f
C1104 a_n10841_1995# dvss 0.502711f
C1105 a_n11219_9395# dvss 0.502711f
C1106 a_n11597_1995# dvss 0.502711f
C1107 a_n11975_9395# dvss 0.502711f
C1108 a_n12353_1995# dvss 0.502711f
C1109 a_n12731_9395# dvss 0.502711f
C1110 a_n13109_1995# dvss 0.502711f
C1111 a_n13487_9395# dvss 0.502711f
C1112 a_n13865_1995# dvss 0.502711f
C1113 a_n14243_9395# dvss 0.502711f
C1114 a_n14621_1995# dvss 0.502711f
C1115 a_n14999_9395# dvss 0.502711f
C1116 dcomp dvss 1.14704f
C1117 comparator_0.n1 dvss 1.33868f
C1118 comparator_0.n0 dvss 0.730766f
C1119 comparator_0.vm dvss 4.47445f
C1120 comparator_0.vn dvss 4.93904f
C1121 ibias_gen_0.ibias dvss 0.498775f
C1122 comparator_0.ena_b dvss 0.625769f
C1123 comparator_0.vnn dvss 22.735302f
C1124 comparator_0.vpp dvss 22.166801f
C1125 ibias_gen_0.ena dvss 5.20891f
C1126 comparator_0.vt dvss 4.0859f
C1127 vl.t0 dvss 6.47511f
C1128 vl.n0 dvss 5.29982f
C1129 sky130_fd_sc_hvl__lsbufhv2lv_1_0.X dvss 0.160791f
C1130 rstring_mux_0.vtrip14.n2 dvss 0.522794f
C1131 rstring_mux_0.vtrip14.n3 dvss 1.031f
C1132 rstring_mux_0.vtrip14.t0 dvss 0.284349f
C1133 rstring_mux_0.vtrip7.n2 dvss 0.400149f
C1134 rstring_mux_0.vtrip7.n3 dvss 1.29459f
C1135 rstring_mux_0.vtrip2.n2 dvss 0.51501f
C1136 rstring_mux_0.vtrip2.n3 dvss 1.03058f
C1137 rstring_mux_0.vtrip2.t4 dvss 0.28851f
C1138 rstring_mux_0.vtrip15.n2 dvss 0.434239f
C1139 rstring_mux_0.vtrip15.n3 dvss 1.28404f
C1140 rstring_mux_0.vtrip3.n2 dvss 0.415891f
C1141 rstring_mux_0.vtrip3.n3 dvss 1.29052f
C1142 rstring_mux_0.vtrip0.n2 dvss 0.523226f
C1143 rstring_mux_0.vtrip0.n3 dvss 1.04554f
C1144 rstring_mux_0.vtrip0.t2 dvss 0.270232f
C1145 rstring_mux_0.vtrip1.n2 dvss 0.423695f
C1146 rstring_mux_0.vtrip1.n3 dvss 1.2886f
C1147 ibias_gen_0.ve.n0 dvss -8.969179f
C1148 ibias_gen_0.ve.t3 dvss 9.08287f
C1149 ibias_gen_0.ve.n2 dvss 0.350991f
C1150 ibias_gen_0.ve.n3 dvss 0.37993f
C1151 ibias_gen_0.ve.n4 dvss 6.82281f
C1152 ibias_gen_0.ve.n5 dvss 7.55903f
C1153 rstring_mux_0.vtrip6.n2 dvss 0.50215f
C1154 rstring_mux_0.vtrip6.n3 dvss 1.02933f
C1155 rstring_mux_0.vtrip6.t2 dvss 0.295855f
C1156 rstring_mux_0.vtop.n0 dvss 0.161879f
C1157 rstring_mux_0.vtop.n1 dvss 0.160951f
C1158 rstring_mux_0.vtop.n2 dvss 0.886062f
C1159 rstring_mux_0.vtop.n3 dvss 0.1411f
C1160 rstring_mux_0.vtop.n4 dvss 0.60016f
C1161 rstring_mux_0.vtop.n5 dvss 0.226235f
C1162 rstring_mux_0.vtop.n6 dvss 0.160951f
C1163 rstring_mux_0.vtop.n7 dvss 0.488298f
C1164 rstring_mux_0.vtop.n8 dvss 0.160951f
C1165 rstring_mux_0.vtop.n9 dvss 0.488298f
C1166 rstring_mux_0.vtop.n10 dvss 0.160951f
C1167 rstring_mux_0.vtop.n11 dvss 0.488298f
C1168 rstring_mux_0.vtop.n12 dvss 0.162293f
C1169 rstring_mux_0.vtop.n13 dvss 0.638369f
C1170 rstring_mux_0.vtop.n14 dvss 0.1411f
C1171 rstring_mux_0.vtop.n15 dvss 0.602669f
C1172 rstring_mux_0.vtop.t0 dvss 4.64098f
C1173 schmitt_trigger_0.in.t7 dvss 2.25707f
C1174 schmitt_trigger_0.in.t14 dvss 1.21543f
C1175 schmitt_trigger_0.in.n5 dvss 1.36804f
C1176 schmitt_trigger_0.in.t12 dvss 1.21543f
C1177 schmitt_trigger_0.in.n6 dvss 1.20717f
C1178 schmitt_trigger_0.in.t6 dvss 1.21543f
C1179 schmitt_trigger_0.in.n7 dvss 1.20717f
C1180 schmitt_trigger_0.in.t13 dvss 1.21543f
C1181 schmitt_trigger_0.in.n8 dvss 1.20717f
C1182 schmitt_trigger_0.in.t9 dvss 1.21543f
C1183 schmitt_trigger_0.in.n9 dvss 1.28817f
C1184 rstring_mux_0.vtrip13.n2 dvss 0.426187f
C1185 rstring_mux_0.vtrip13.n3 dvss 1.28724f
C1186 rstring_mux_0.vtrip4.n2 dvss 0.508844f
C1187 rstring_mux_0.vtrip4.n3 dvss 1.02973f
C1188 rstring_mux_0.vtrip4.t0 dvss 0.292274f
C1189 rstring_mux_0.vtrip5.n2 dvss 0.405641f
C1190 rstring_mux_0.vtrip5.n3 dvss 1.29292f
C1191 ibias_gen_0.vstart.n0 dvss 1.41043f
C1192 ibias_gen_0.vstart.n1 dvss 0.258324f
C1193 ibias_gen_0.vstart.t0 dvss 0.344828f
C1194 ibias_gen_0.vstart.n2 dvss 0.255572f
C1195 ibias_gen_0.vstart.n3 dvss 0.260069f
C1196 ibias_gen_0.vstart.n4 dvss 0.255572f
C1197 ibias_gen_0.vstart.n5 dvss 0.750761f
C1198 ibias_gen_0.vstart.n6 dvss 0.398642f
C1199 ibias_gen_0.vstart.n7 dvss 0.255572f
C1200 rstring_mux_0.vtrip11.n2 dvss 0.418122f
C1201 rstring_mux_0.vtrip11.n3 dvss 1.28961f
C1202 vbg_1v2.t24 dvss 1.08995f
C1203 vbg_1v2.t2 dvss 1.07574f
C1204 vbg_1v2.n0 dvss 0.859433f
C1205 vbg_1v2.t0 dvss 1.07574f
C1206 vbg_1v2.n1 dvss 0.44661f
C1207 vbg_1v2.t4 dvss 1.07574f
C1208 vbg_1v2.n2 dvss 0.44661f
C1209 vbg_1v2.t7 dvss 1.07574f
C1210 vbg_1v2.n3 dvss 0.44661f
C1211 vbg_1v2.t6 dvss 1.07574f
C1212 vbg_1v2.n4 dvss 0.44661f
C1213 vbg_1v2.t11 dvss 1.07574f
C1214 vbg_1v2.n5 dvss 0.44661f
C1215 vbg_1v2.t9 dvss 1.07574f
C1216 vbg_1v2.n6 dvss 0.665796f
C1217 vbg_1v2.t8 dvss 1.10059f
C1218 vbg_1v2.t14 dvss 1.08611f
C1219 vbg_1v2.n7 dvss 0.883289f
C1220 vbg_1v2.t13 dvss 1.08611f
C1221 vbg_1v2.n8 dvss 0.458671f
C1222 vbg_1v2.t17 dvss 1.08611f
C1223 vbg_1v2.n9 dvss 0.458671f
C1224 vbg_1v2.t20 dvss 1.08611f
C1225 vbg_1v2.n10 dvss 0.458671f
C1226 vbg_1v2.t18 dvss 1.08611f
C1227 vbg_1v2.n11 dvss 0.458671f
C1228 vbg_1v2.t23 dvss 1.08611f
C1229 vbg_1v2.n12 dvss 0.458671f
C1230 vbg_1v2.t21 dvss 1.08611f
C1231 vbg_1v2.n13 dvss 0.608433f
C1232 vbg_1v2.n14 dvss 1.8485f
C1233 vbg_1v2.n15 dvss 0.183619f
C1234 vbg_1v2.n16 dvss 0.144543f
C1235 vbg_1v2.n17 dvss 0.144543f
C1236 vbg_1v2.n18 dvss 0.144543f
C1237 vbg_1v2.n19 dvss 0.282418f
C1238 vbg_1v2.t22 dvss 0.419943f
C1239 vbg_1v2.t19 dvss 0.419596f
C1240 vbg_1v2.n20 dvss 0.282418f
C1241 vbg_1v2.n21 dvss 0.144543f
C1242 vbg_1v2.t15 dvss 0.419596f
C1243 vbg_1v2.n22 dvss 0.144543f
C1244 vbg_1v2.t12 dvss 0.419596f
C1245 vbg_1v2.n23 dvss 0.144543f
C1246 vbg_1v2.n24 dvss 0.144543f
C1247 vbg_1v2.t5 dvss 0.419596f
C1248 vbg_1v2.n25 dvss 0.144543f
C1249 vbg_1v2.t3 dvss 0.419596f
C1250 vbg_1v2.n26 dvss 0.144543f
C1251 vbg_1v2.n27 dvss 0.144543f
C1252 vbg_1v2.t1 dvss 0.419596f
C1253 vbg_1v2.n28 dvss 0.144543f
C1254 vbg_1v2.t25 dvss 0.419596f
C1255 vbg_1v2.n29 dvss 0.144543f
C1256 vbg_1v2.n30 dvss 0.143946f
C1257 vbg_1v2.t10 dvss 0.419596f
C1258 vbg_1v2.n31 dvss 0.143946f
C1259 vbg_1v2.t16 dvss 0.419596f
C1260 vbg_1v2.n32 dvss 0.134129f
C1261 vbg_1v2.n33 dvss 0.213865f
C1262 ibias_gen_0.vn1.n0 dvss 0.762542f
C1263 ibias_gen_0.vn1.t4 dvss 2.16042f
C1264 ibias_gen_0.vn1.t15 dvss 2.16042f
C1265 ibias_gen_0.vn1.t10 dvss 2.24798f
C1266 ibias_gen_0.vn1.n2 dvss 1.43288f
C1267 ibias_gen_0.vn1.t17 dvss 2.16042f
C1268 ibias_gen_0.vn1.t14 dvss 2.24798f
C1269 ibias_gen_0.vn1.n3 dvss 1.40011f
C1270 ibias_gen_0.vn1.n4 dvss 0.14406f
C1271 ibias_gen_0.vn1.t11 dvss 2.16042f
C1272 ibias_gen_0.vn1.t12 dvss 2.24798f
C1273 ibias_gen_0.vn1.n5 dvss 1.43288f
C1274 ibias_gen_0.vn1.t13 dvss 2.16042f
C1275 ibias_gen_0.vn1.t16 dvss 2.24798f
C1276 ibias_gen_0.vn1.n6 dvss 1.40011f
C1277 ibias_gen_0.vn1.n7 dvss 0.14406f
C1278 ibias_gen_0.vn1.n8 dvss 0.113548f
C1279 ibias_gen_0.vn1.n9 dvss 0.721953f
C1280 ibias_gen_0.vn1.t6 dvss 2.20687f
C1281 ibias_gen_0.vn1.n10 dvss 0.735436f
C1282 ibias_gen_0.vn1.n12 dvss 0.223089f
C1283 ibias_gen_0.vn1.n13 dvss 0.123215f
C1284 ibias_gen_0.vp1.n0 dvss 2.00743f
C1285 ibias_gen_0.vp1.t13 dvss 2.42566f
C1286 ibias_gen_0.vp1.n1 dvss 0.11654f
C1287 ibias_gen_0.vp1.n2 dvss 0.22885f
C1288 ibias_gen_0.vp1.n3 dvss 1.906f
C1289 ibias_gen_0.vp1.t15 dvss 2.42228f
C1290 ibias_gen_0.vp1.n4 dvss 0.20081f
C1291 ibias_gen_0.vp1.n5 dvss 0.870858f
C1292 ibias_gen_0.vp1.n6 dvss 0.137903f
C1293 ibias_gen_0.vp1.n7 dvss 0.190001f
C1294 ibias_gen_0.vp1.n8 dvss 0.150339f
C1295 ibias_gen_0.vp1.n9 dvss 0.888932f
C1296 ibias_gen_0.vp1.n10 dvss 0.150339f
C1297 ibias_gen_0.vp1.n11 dvss 0.603419f
C1298 ibias_gen_0.vp1.n12 dvss 0.145319f
C1299 ibias_gen_0.vp1.n13 dvss 0.592886f
C1300 ibias_gen_0.vp1.n14 dvss 0.176014f
C1301 ibias_gen_0.vp1.n15 dvss 0.738575f
C1302 schmitt_trigger_0.m.n3 dvss 0.65613f
C1303 schmitt_trigger_0.m.n4 dvss 0.195435f
C1304 schmitt_trigger_0.m.n7 dvss 0.732652f
C1305 schmitt_trigger_0.m.t17 dvss 0.161114f
C1306 schmitt_trigger_0.m.t14 dvss 0.164304f
C1307 schmitt_trigger_0.m.t15 dvss 0.16415f
C1308 schmitt_trigger_0.m.n8 dvss 0.16975f
C1309 schmitt_trigger_0.m.t16 dvss 0.16428f
C1310 schmitt_trigger_0.m.n9 dvss 0.374799f
C1311 schmitt_trigger_0.m.n10 dvss 0.537335f
C1312 schmitt_trigger_0.m.n11 dvss 0.312554f
C1313 schmitt_trigger_0.m.n13 dvss 0.192206f
C1314 schmitt_trigger_0.m.n15 dvss 0.222965f
C1315 rstring_mux_0.vtrip10.n2 dvss 0.511346f
C1316 rstring_mux_0.vtrip10.n3 dvss 1.02889f
C1317 rstring_mux_0.vtrip10.t2 dvss 0.291299f
C1318 ibias_gen_0.vp.n0 dvss 0.409208f
C1319 ibias_gen_0.vp.t4 dvss 0.178419f
C1320 ibias_gen_0.vp.n3 dvss 0.627732f
C1321 ibias_gen_0.vp.t10 dvss 1.62254f
C1322 ibias_gen_0.vp.n4 dvss 1.22303f
C1323 ibias_gen_0.vp.t8 dvss 1.56547f
C1324 ibias_gen_0.vp.n5 dvss 1.22303f
C1325 ibias_gen_0.vp.t7 dvss 1.56547f
C1326 ibias_gen_0.vp.n6 dvss 1.22303f
C1327 ibias_gen_0.vp.t9 dvss 1.594f
C1328 ibias_gen_0.vp.n7 dvss 0.744925f
C1329 ibias_gen_0.vp.n8 dvss 0.92267f
C1330 ibias_gen_0.vp.n10 dvss 0.463021f
C1331 ibias_gen_0.vr.n0 dvss 0.183081f
C1332 ibias_gen_0.vr.n1 dvss 0.161866f
C1333 ibias_gen_0.vr.n2 dvss 1.54735f
C1334 ibias_gen_0.vr.t4 dvss 0.540543f
C1335 ibias_gen_0.vp0.n0 dvss 0.799876f
C1336 ibias_gen_0.vp0.n1 dvss 0.223451f
C1337 ibias_gen_0.vp0.n3 dvss 0.912302f
C1338 ibias_gen_0.vp0.n5 dvss 0.161869f
C1339 ibias_gen_0.vp0.t2 dvss 1.77926f
C1340 ibias_gen_0.vp0.n6 dvss 1.51784f
C1341 ibias_gen_0.vp0.n7 dvss 0.745969f
C1342 ibias_gen_0.vp0.t13 dvss 1.81292f
C1343 ibias_gen_0.vp0.t12 dvss 1.74916f
C1344 ibias_gen_0.vp0.n8 dvss 1.51784f
C1345 ibias_gen_0.vp0.n9 dvss 0.824132f
C1346 ibias_gen_0.vp0.t4 dvss 1.74916f
C1347 ibias_gen_0.vp0.n10 dvss 0.822001f
C1348 ibias_gen_0.vp0.n11 dvss 0.13184f
C1349 ibias_gen_0.vp0.n12 dvss 1.01161f
C1350 ibias_gen_0.vp0.n13 dvss 1.10668f
C1351 ibias_gen_0.vp0.n14 dvss 0.143186f
C1352 ibias_gen_0.Mt4 dvss 1.25878f
C1353 ibias_gen_0.vn0.n0 dvss 0.935654f
C1354 ibias_gen_0.vn0.n1 dvss 1.39652f
C1355 ibias_gen_0.vn0.n2 dvss 0.142325f
C1356 ibias_gen_0.vn0.n3 dvss 0.874872f
C1357 ibias_gen_0.vn0.t19 dvss 2.24075f
C1358 ibias_gen_0.vn0.t3 dvss 2.19836f
C1359 ibias_gen_0.vn0.n4 dvss 0.920525f
C1360 ibias_gen_0.vn0.n5 dvss 0.111014f
C1361 ibias_gen_0.vn0.n6 dvss 0.198283f
C1362 ibias_gen_0.vn0.n7 dvss 0.161371f
C1363 ibias_gen_0.vn0.t1 dvss 2.16084f
C1364 ibias_gen_0.vn0.n8 dvss 1.01955f
C1365 ibias_gen_0.vn0.n9 dvss 1.87632f
C1366 ibias_gen_0.vn0.t20 dvss 2.16084f
C1367 ibias_gen_0.vn0.n10 dvss 1.71213f
C1368 ibias_gen_0.vn0.n11 dvss 0.975041f
C1369 ibias_gen_0.vn0.t13 dvss 0.202556f
C1370 ibias_gen_0.vn0.n12 dvss 0.12274f
C1371 ibias_gen_0.vn0.n13 dvss 0.12274f
C1372 ibias_gen_0.vn0.n14 dvss 0.12274f
C1373 ibias_gen_0.vn0.n15 dvss 0.12274f
C1374 ibias_gen_0.vn0.n16 dvss 0.12274f
C1375 dvdd.t4 dvss 0.108773f
C1376 dvdd.t125 dvss 0.108773f
C1377 dvdd.t138 dvss 0.108773f
C1378 dvdd.t100 dvss 0.108773f
C1379 dvdd.t94 dvss 0.108773f
C1380 dvdd.t92 dvss 0.108773f
C1381 dvdd.t116 dvss 0.108773f
C1382 dvdd.t80 dvss 0.108773f
C1383 dvdd.t96 dvss 0.108773f
C1384 dvdd.n99 dvss 0.135907f
C1385 dvdd.n105 dvss 0.127548f
C1386 dvdd.n117 dvss 0.233166f
C1387 dvdd.t102 dvss 0.212041f
C1388 dvdd.t104 dvss 0.172483f
C1389 dvdd.t106 dvss 0.172483f
C1390 dvdd.t121 dvss 0.172483f
C1391 dvdd.t68 dvss 0.172483f
C1392 dvdd.t64 dvss 0.172483f
C1393 dvdd.t60 dvss 0.172483f
C1394 dvdd.t16 dvss 0.172483f
C1395 dvdd.t18 dvss 0.172483f
C1396 dvdd.t24 dvss 0.172483f
C1397 dvdd.t14 dvss 0.172483f
C1398 dvdd.t20 dvss 0.172483f
C1399 dvdd.t22 dvss 0.212041f
C1400 dvdd.n118 dvss 0.233166f
C1401 dvdd.n121 dvss 0.104808f
C1402 dvdd.n122 dvss 0.309736f
C1403 dvdd.t42 dvss 0.133335f
C1404 dvdd.n179 dvss 0.180651f
C1405 dvdd.n180 dvss 0.332137f
C1406 dvdd.n181 dvss 0.722016f
C1407 dvdd.n182 dvss 0.722016f
C1408 dvdd.n183 dvss 2.69721f
C1409 dvdd.n184 dvss 0.332827f
C1410 dvdd.n185 dvss 0.725257f
C1411 dvdd.n186 dvss 2.7446f
C1412 dvdd.n187 dvss 2.69721f
C1413 dvdd.n188 dvss 2.7446f
C1414 dvdd.n189 dvss 0.725257f
C1415 dvdd.n190 dvss 0.316688f
C1416 dvdd.n191 dvss 0.176035f
C1417 dvdd.n193 dvss 1.47224f
C1418 dvdd.t12 dvss 0.108773f
C1419 dvdd.t127 dvss 0.108773f
C1420 dvdd.t129 dvss 0.108773f
C1421 dvdd.t114 dvss 0.108773f
C1422 dvdd.t0 dvss 0.108773f
C1423 dvdd.t86 dvss 0.108773f
C1424 dvdd.t123 dvss 0.108773f
C1425 dvdd.t98 dvss 0.108773f
C1426 dvdd.t2 dvss 0.108773f
C1427 dvdd.t112 dvss 0.150767f
C1428 dvdd.t131 dvss 0.141125f
C1429 dvdd.n302 dvss 1.29926f
C1430 dvdd.n303 dvss 1.16605f
C1431 schmitt_trigger_0.out.n5 dvss 0.689226f
C1432 schmitt_trigger_0.out.t6 dvss 0.155689f
C1433 schmitt_trigger_0.out.t12 dvss 0.155538f
C1434 schmitt_trigger_0.out.n6 dvss 0.163942f
C1435 schmitt_trigger_0.out.t15 dvss 0.155622f
C1436 schmitt_trigger_0.out.n7 dvss 0.113412f
C1437 schmitt_trigger_0.out.t8 dvss 0.162392f
C1438 schmitt_trigger_0.out.n8 dvss 0.688643f
C1439 schmitt_trigger_0.out.n9 dvss 0.41845f
C1440 schmitt_trigger_0.out.n10 dvss 0.606738f
C1441 schmitt_trigger_0.out.n11 dvss 0.342028f
C1442 rstring_mux_0.vtrip8.n2 dvss 0.503767f
C1443 rstring_mux_0.vtrip8.n3 dvss 1.02946f
C1444 rstring_mux_0.vtrip8.t2 dvss 0.294942f
C1445 rstring_mux_0.vtrip9.n2 dvss 0.409678f
C1446 rstring_mux_0.vtrip9.n3 dvss 1.29226f
C1447 avdd.t206 dvss 2.41161f
C1448 avdd.t381 dvss 0.98697f
C1449 avdd.t328 dvss 1.6121f
C1450 avdd.t181 dvss 2.41161f
C1451 avdd.t325 dvss 0.98697f
C1452 avdd.t189 dvss 1.6121f
C1453 avdd.t214 dvss 2.41161f
C1454 avdd.t351 dvss 0.98697f
C1455 avdd.t10 dvss 1.6121f
C1456 avdd.t284 dvss 2.41161f
C1457 avdd.t373 dvss 0.98697f
C1458 avdd.t330 dvss 1.6121f
C1459 avdd.t274 dvss 2.41161f
C1460 avdd.t272 dvss 0.98697f
C1461 avdd.t282 dvss 1.6121f
C1462 avdd.t318 dvss 2.41161f
C1463 avdd.t316 dvss 0.98697f
C1464 avdd.t253 dvss 1.6121f
C1465 avdd.t187 dvss 2.41161f
C1466 avdd.t286 dvss 0.98697f
C1467 avdd.t248 dvss 1.6121f
C1468 avdd.t379 dvss 2.41161f
C1469 avdd.t377 dvss 0.98697f
C1470 avdd.t303 dvss 1.6121f
C1471 avdd.t360 dvss 0.323361f
C1472 avdd.n69 dvss 0.785005f
C1473 avdd.n73 dvss 0.177625f
C1474 avdd.n74 dvss 0.794328f
C1475 avdd.n75 dvss 2.86889f
C1476 avdd.t296 dvss 1.69812f
C1477 avdd.n78 dvss 1.28424f
C1478 avdd.n83 dvss 0.102203f
C1479 avdd.n88 dvss 0.271799f
C1480 avdd.n90 dvss 0.10665f
C1481 avdd.n94 dvss 0.609671f
C1482 avdd.t354 dvss 0.323361f
C1483 avdd.n95 dvss 0.360413f
C1484 avdd.n96 dvss 0.518725f
C1485 avdd.n99 dvss 0.451358f
C1486 avdd.n100 dvss 0.646723f
C1487 avdd.t358 dvss 1.58312f
C1488 avdd.t260 dvss 0.289678f
C1489 avdd.n101 dvss 0.586092f
C1490 avdd.n116 dvss 0.102203f
C1491 avdd.n119 dvss 0.271799f
C1492 avdd.n124 dvss 0.10665f
C1493 avdd.n126 dvss 1.69528f
C1494 avdd.n129 dvss 1.43803f
C1495 avdd.n144 dvss 0.102203f
C1496 avdd.n147 dvss 0.271799f
C1497 avdd.n152 dvss 0.10665f
C1498 avdd.n154 dvss 1.69528f
C1499 avdd.n157 dvss 1.43803f
C1500 avdd.n172 dvss 0.102203f
C1501 avdd.n175 dvss 0.271799f
C1502 avdd.n180 dvss 0.10665f
C1503 avdd.n182 dvss 1.69528f
C1504 avdd.n185 dvss 1.43803f
C1505 avdd.n200 dvss 0.102203f
C1506 avdd.n203 dvss 0.271799f
C1507 avdd.n208 dvss 0.10665f
C1508 avdd.n210 dvss 1.69528f
C1509 avdd.n213 dvss 1.43803f
C1510 avdd.n228 dvss 0.102203f
C1511 avdd.n231 dvss 0.271799f
C1512 avdd.n236 dvss 0.10665f
C1513 avdd.n238 dvss 1.69528f
C1514 avdd.n241 dvss 1.43803f
C1515 avdd.n256 dvss 0.102203f
C1516 avdd.n259 dvss 0.271799f
C1517 avdd.n264 dvss 0.10665f
C1518 avdd.n266 dvss 1.69528f
C1519 avdd.n269 dvss 1.43803f
C1520 avdd.n284 dvss 0.102203f
C1521 avdd.n287 dvss 0.271799f
C1522 avdd.n292 dvss 0.10665f
C1523 avdd.n294 dvss 1.69528f
C1524 avdd.n297 dvss 1.43803f
C1525 avdd.n312 dvss 0.102203f
C1526 avdd.n315 dvss 0.271799f
C1527 avdd.n320 dvss 0.10665f
C1528 avdd.n322 dvss 1.69528f
C1529 avdd.n325 dvss 1.43803f
C1530 avdd.t268 dvss 2.41161f
C1531 avdd.t313 dvss 0.98697f
C1532 avdd.t276 dvss 1.6121f
C1533 avdd.t8 dvss 2.41161f
C1534 avdd.t6 dvss 0.98697f
C1535 avdd.t191 dvss 1.6121f
C1536 avdd.t2 dvss 2.41161f
C1537 avdd.t0 dvss 0.98697f
C1538 avdd.t305 dvss 1.6121f
C1539 avdd.t70 dvss 2.41161f
C1540 avdd.t74 dvss 0.98697f
C1541 avdd.t294 dvss 1.6121f
C1542 avdd.t193 dvss 2.41161f
C1543 avdd.t195 dvss 0.98697f
C1544 avdd.t183 dvss 1.6121f
C1545 avdd.t280 dvss 2.41161f
C1546 avdd.t290 dvss 0.98697f
C1547 avdd.t370 dvss 1.6121f
C1548 avdd.t208 dvss 2.41161f
C1549 avdd.t258 dvss 0.98697f
C1550 avdd.t292 dvss 1.6121f
C1551 avdd.t72 dvss 2.41161f
C1552 avdd.t251 dvss 0.98697f
C1553 avdd.t307 dvss 1.6121f
C1554 avdd.t242 dvss 2.18605f
C1555 avdd.t240 dvss 0.894656f
C1556 avdd.t255 dvss 1.52814f
C1557 avdd.n408 dvss 1.86981f
C1558 avdd.n409 dvss 0.102203f
C1559 avdd.n417 dvss 0.271799f
C1560 avdd.n419 dvss 0.10665f
C1561 avdd.n423 dvss 1.30352f
C1562 avdd.n438 dvss 0.102203f
C1563 avdd.n441 dvss 0.271799f
C1564 avdd.n446 dvss 0.10665f
C1565 avdd.n448 dvss 1.69528f
C1566 avdd.n451 dvss 1.43803f
C1567 avdd.n466 dvss 0.102203f
C1568 avdd.n469 dvss 0.271799f
C1569 avdd.n474 dvss 0.10665f
C1570 avdd.n476 dvss 1.69528f
C1571 avdd.n479 dvss 1.43803f
C1572 avdd.n494 dvss 0.102203f
C1573 avdd.n497 dvss 0.271799f
C1574 avdd.n502 dvss 0.10665f
C1575 avdd.n504 dvss 1.69528f
C1576 avdd.n507 dvss 1.43803f
C1577 avdd.n522 dvss 0.102203f
C1578 avdd.n525 dvss 0.271799f
C1579 avdd.n530 dvss 0.10665f
C1580 avdd.n532 dvss 1.69528f
C1581 avdd.n535 dvss 1.43803f
C1582 avdd.n550 dvss 0.102203f
C1583 avdd.n553 dvss 0.271799f
C1584 avdd.n558 dvss 0.10665f
C1585 avdd.n560 dvss 1.69528f
C1586 avdd.n563 dvss 1.43803f
C1587 avdd.n578 dvss 0.102203f
C1588 avdd.n581 dvss 0.271799f
C1589 avdd.n586 dvss 0.10665f
C1590 avdd.n588 dvss 1.69528f
C1591 avdd.n591 dvss 1.43803f
C1592 avdd.n606 dvss 0.102203f
C1593 avdd.n609 dvss 0.271799f
C1594 avdd.n614 dvss 0.10665f
C1595 avdd.n616 dvss 1.69528f
C1596 avdd.n619 dvss 1.43803f
C1597 avdd.n634 dvss 0.102203f
C1598 avdd.n637 dvss 0.271799f
C1599 avdd.n642 dvss 0.10665f
C1600 avdd.n644 dvss 1.69528f
C1601 avdd.n647 dvss 1.43803f
C1602 avdd.n659 dvss 5.72462f
C1603 avdd.n660 dvss 7.31017f
C1604 avdd.n661 dvss 6.43982f
C1605 avdd.t333 dvss 0.111115f
C1606 avdd.t332 dvss 1.21874f
C1607 avdd.n667 dvss 0.722284f
C1608 avdd.n673 dvss 0.372238f
C1609 avdd.n674 dvss 0.140742f
C1610 avdd.n675 dvss 1.32173f
C1611 avdd.t91 dvss 0.947086f
C1612 avdd.n676 dvss 0.588009f
C1613 avdd.n677 dvss 1.29698f
C1614 avdd.n678 dvss 0.775203f
C1615 avdd.n679 dvss 2.55802f
C1616 avdd.n680 dvss 2.55802f
C1617 avdd.n681 dvss 0.775203f
C1618 avdd.n682 dvss 1.29759f
C1619 avdd.n684 dvss 0.384107f
C1620 avdd.t185 dvss 0.60848f
C1621 avdd.n691 dvss 0.228763f
C1622 avdd.n692 dvss 1.0121f
C1623 avdd.n693 dvss 1.00517f
C1624 avdd.t429 dvss 0.221831f
C1625 avdd.t270 dvss 0.221831f
C1626 avdd.t430 dvss 0.111115f
C1627 avdd.n702 dvss 0.372238f
C1628 avdd.n704 dvss 0.256492f
C1629 avdd.n710 dvss 0.228763f
C1630 avdd.n712 dvss 1.0121f
C1631 avdd.n713 dvss 1.00517f
C1632 avdd.t38 dvss 0.221831f
C1633 avdd.t264 dvss 0.221831f
C1634 avdd.t39 dvss 0.111115f
C1635 avdd.n722 dvss 0.372238f
C1636 avdd.n724 dvss 0.256492f
C1637 avdd.n730 dvss 0.228763f
C1638 avdd.n732 dvss 1.0121f
C1639 avdd.n733 dvss 1.00517f
C1640 avdd.t299 dvss 0.221831f
C1641 avdd.t216 dvss 0.221831f
C1642 avdd.t300 dvss 0.111115f
C1643 avdd.n742 dvss 0.372238f
C1644 avdd.n744 dvss 0.256492f
C1645 avdd.n750 dvss 0.228763f
C1646 avdd.n752 dvss 1.0121f
C1647 avdd.n753 dvss 1.00517f
C1648 avdd.t68 dvss 0.221831f
C1649 avdd.t36 dvss 0.221831f
C1650 avdd.t69 dvss 0.111115f
C1651 avdd.n762 dvss 0.372238f
C1652 avdd.n764 dvss 0.256492f
C1653 avdd.n770 dvss 0.228763f
C1654 avdd.n772 dvss 1.0121f
C1655 avdd.n773 dvss 1.00517f
C1656 avdd.t437 dvss 0.221831f
C1657 avdd.t419 dvss 0.794121f
C1658 avdd.t438 dvss 0.111115f
C1659 avdd.n782 dvss 0.372238f
C1660 avdd.n784 dvss 0.256492f
C1661 avdd.n785 dvss 0.2691f
C1662 avdd.n786 dvss 0.19407f
C1663 avdd.t420 dvss 0.111115f
C1664 avdd.n789 dvss 0.372238f
C1665 avdd.n795 dvss 1.00517f
C1666 avdd.n796 dvss 1.0121f
C1667 avdd.n797 dvss 0.228763f
C1668 avdd.n801 dvss 0.256492f
C1669 avdd.t279 dvss 0.111115f
C1670 avdd.n802 dvss 0.372238f
C1671 avdd.n807 dvss 1.0121f
C1672 avdd.n808 dvss 0.228763f
C1673 avdd.t278 dvss 0.221831f
C1674 avdd.n809 dvss 1.00517f
C1675 avdd.n812 dvss 0.256492f
C1676 avdd.t37 dvss 0.111115f
C1677 avdd.n814 dvss 0.372238f
C1678 avdd.n820 dvss 1.00517f
C1679 avdd.n821 dvss 1.0121f
C1680 avdd.n822 dvss 0.228763f
C1681 avdd.n826 dvss 0.256492f
C1682 avdd.t239 dvss 0.111115f
C1683 avdd.n827 dvss 0.372238f
C1684 avdd.n832 dvss 1.0121f
C1685 avdd.n833 dvss 0.228763f
C1686 avdd.t238 dvss 0.221831f
C1687 avdd.n834 dvss 1.00517f
C1688 avdd.n837 dvss 0.256492f
C1689 avdd.t217 dvss 0.111115f
C1690 avdd.n839 dvss 0.372238f
C1691 avdd.n845 dvss 1.00517f
C1692 avdd.n846 dvss 1.0121f
C1693 avdd.n847 dvss 0.228763f
C1694 avdd.n851 dvss 0.256492f
C1695 avdd.t198 dvss 0.111115f
C1696 avdd.n852 dvss 0.372238f
C1697 avdd.n857 dvss 1.0121f
C1698 avdd.n858 dvss 0.228763f
C1699 avdd.t197 dvss 0.221831f
C1700 avdd.n859 dvss 1.00517f
C1701 avdd.n862 dvss 0.256492f
C1702 avdd.t265 dvss 0.111115f
C1703 avdd.n864 dvss 0.372238f
C1704 avdd.n870 dvss 1.00517f
C1705 avdd.n871 dvss 1.0121f
C1706 avdd.n872 dvss 0.228763f
C1707 avdd.n876 dvss 0.256492f
C1708 avdd.t432 dvss 0.111115f
C1709 avdd.n877 dvss 0.372238f
C1710 avdd.n882 dvss 1.0121f
C1711 avdd.n883 dvss 0.228763f
C1712 avdd.t431 dvss 0.221831f
C1713 avdd.n884 dvss 1.00517f
C1714 avdd.n887 dvss 0.256492f
C1715 avdd.t271 dvss 0.111115f
C1716 avdd.n889 dvss 0.372238f
C1717 avdd.n895 dvss 1.00517f
C1718 avdd.n896 dvss 1.0121f
C1719 avdd.n897 dvss 0.228763f
C1720 avdd.n901 dvss 0.256492f
C1721 avdd.t267 dvss 0.111115f
C1722 avdd.n902 dvss 0.372238f
C1723 avdd.n907 dvss 1.0121f
C1724 avdd.n908 dvss 0.228763f
C1725 avdd.t266 dvss 0.221831f
C1726 avdd.n909 dvss 1.00517f
C1727 avdd.n912 dvss 0.256492f
C1728 avdd.t186 dvss 0.111115f
C1729 avdd.n913 dvss 0.372238f
C1730 avdd.n919 dvss 1.25828f
C1731 avdd.t126 dvss 0.947086f
C1732 avdd.t89 dvss 0.947086f
C1733 avdd.t139 dvss 0.947086f
C1734 avdd.t111 dvss 0.947086f
C1735 avdd.t162 dvss 0.947086f
C1736 avdd.t102 dvss 0.947086f
C1737 avdd.t177 dvss 0.947086f
C1738 avdd.t166 dvss 0.947086f
C1739 avdd.t156 dvss 0.947086f
C1740 avdd.t164 dvss 0.947086f
C1741 avdd.t124 dvss 0.947086f
C1742 avdd.t175 dvss 0.947086f
C1743 avdd.t179 dvss 0.947086f
C1744 avdd.t151 dvss 0.947086f
C1745 avdd.n920 dvss 0.589555f
C1746 avdd.n921 dvss 0.589555f
C1747 avdd.n922 dvss 0.589555f
C1748 avdd.n923 dvss 0.589555f
C1749 avdd.n924 dvss 0.589555f
C1750 avdd.n925 dvss 0.589555f
C1751 avdd.n926 dvss 0.460172f
C1752 avdd.n927 dvss 0.137631f
C1753 avdd.n928 dvss 0.581308f
C1754 avdd.n929 dvss 0.589555f
C1755 avdd.n930 dvss 0.589555f
C1756 avdd.n931 dvss 0.589555f
C1757 avdd.n932 dvss 0.589555f
C1758 avdd.n933 dvss 0.589555f
C1759 avdd.n934 dvss 0.605506f
C1760 avdd.n935 dvss 0.374869f
C1761 avdd.n936 dvss 3.03751f
C1762 avdd.n937 dvss 11.6733f
C1763 avdd.n938 dvss 1.00206f
C1764 avdd.n939 dvss 3.2921f
C1765 avdd.t133 dvss 2.10465f
C1766 avdd.n940 dvss 1.34047f
C1767 avdd.n941 dvss 0.120301f
C1768 avdd.n942 dvss 1.4146f
C1769 avdd.n943 dvss 0.948991f
C1770 avdd.n944 dvss 0.221947f
C1771 avdd.n945 dvss 0.174834f
C1772 avdd.n946 dvss 0.240832f
C1773 avdd.n947 dvss 0.322853f
C1774 avdd.n948 dvss 0.547718f
C1775 avdd.n949 dvss 0.547718f
C1776 avdd.t342 dvss 1.85494f
C1777 avdd.t80 dvss 36.501698f
C1778 avdd.n950 dvss 1.45348f
C1779 avdd.n951 dvss 3.24482f
C1780 avdd.n952 dvss 1.6959f
C1781 avdd.n953 dvss 1.03094f
C1782 avdd.t14 dvss 34.6356f
C1783 avdd.t17 dvss 46.1808f
C1784 avdd.t21 dvss 34.6356f
C1785 avdd.n954 dvss 1.45348f
C1786 avdd.n955 dvss 0.869726f
C1787 avdd.n956 dvss 0.869726f
C1788 avdd.n957 dvss 1.90685f
C1789 avdd.n958 dvss 1.4146f
C1790 avdd.n960 dvss 0.29269f
C1791 avdd.n961 dvss 1.4854f
C1792 avdd.n962 dvss 1.96715f
C1793 avdd.n963 dvss 1.93091f
C1794 avdd.n964 dvss 1.12799f
C1795 avdd.n965 dvss 1.07468f
C1796 avdd.n966 dvss 0.140283f
C1797 avdd.n967 dvss 0.140209f
C1798 avdd.n968 dvss 1.01373f
C1799 avdd.n969 dvss 1.4146f
C1800 avdd.n970 dvss 0.294294f
C1801 avdd.n971 dvss 0.352378f
C1802 avdd.n972 dvss 0.387122f
C1803 avdd.n973 dvss 0.656852f
C1804 avdd.n974 dvss 0.656852f
C1805 avdd.t12 dvss 46.1808f
C1806 avdd.t84 dvss 36.501698f
C1807 avdd.n975 dvss 1.93486f
C1808 avdd.n976 dvss 14.734401f
C1809 avdd.n978 dvss 0.347625f
C1810 avdd.n980 dvss 0.347625f
C1811 avdd.n982 dvss 0.347625f
C1812 avdd.n984 dvss 0.347625f
C1813 avdd.n985 dvss 0.373633f
C1814 avdd.n986 dvss 0.230478f
C1815 avdd.n987 dvss 0.210423f
C1816 avdd.n988 dvss 1.87616f
C1817 avdd.t246 dvss 1.41679f
C1818 avdd.t244 dvss 1.14534f
C1819 avdd.t54 dvss 1.14534f
C1820 avdd.t64 dvss 1.14534f
C1821 avdd.t62 dvss 0.859008f
C1822 avdd.n989 dvss 1.8957f
C1823 avdd.t58 dvss 0.859008f
C1824 avdd.t66 dvss 1.14534f
C1825 avdd.t60 dvss 1.14534f
C1826 avdd.t56 dvss 1.14534f
C1827 avdd.t52 dvss 1.41679f
C1828 avdd.n990 dvss 1.87616f
C1829 avdd.n991 dvss 0.210423f
C1830 avdd.n992 dvss 0.228974f
C1831 avdd.n993 dvss 0.298278f
C1832 avdd.n994 dvss 2.05986f
C1833 avdd.n995 dvss 0.141631f
C1834 avdd.n996 dvss 0.140283f
C1835 avdd.n998 dvss 0.195382f
C1836 avdd.n1000 dvss 0.196804f
C1837 avdd.n1002 dvss 0.196804f
C1838 avdd.n1004 dvss 0.196804f
C1839 avdd.n1006 dvss 0.196804f
C1840 avdd.n1008 dvss 0.196804f
C1841 avdd.n1010 dvss 0.196804f
C1842 avdd.n1012 dvss 0.196804f
C1843 avdd.n1014 dvss 0.175474f
C1844 avdd.t344 dvss 2.04059f
C1845 avdd.n1015 dvss 1.75782f
C1846 avdd.n1016 dvss 0.20375f
C1847 avdd.n1017 dvss 0.188858f
C1848 avdd.n1018 dvss 1.01121f
C1849 avdd.n1019 dvss 1.75491f
C1850 avdd.n1020 dvss 1.88613f
C1851 avdd.n1021 dvss 0.257938f
C1852 avdd.n1022 dvss 4.38252f
C1853 avdd.n1023 dvss 3.2921f
C1854 avdd.n1024 dvss 0.257938f
C1855 avdd.n1025 dvss 0.196804f
C1856 avdd.t83 dvss 2.10465f
C1857 avdd.n1026 dvss 0.141631f
C1858 avdd.t104 dvss 2.10465f
C1859 avdd.n1027 dvss 1.34047f
C1860 avdd.n1029 dvss 0.195382f
C1861 avdd.n1030 dvss 0.196804f
C1862 avdd.t116 dvss 2.10465f
C1863 avdd.t173 dvss 2.10465f
C1864 avdd.n1032 dvss 1.34047f
C1865 avdd.n1033 dvss 0.141631f
C1866 avdd.n1034 dvss 0.141631f
C1867 avdd.n1035 dvss 1.34047f
C1868 avdd.n1037 dvss 0.196804f
C1869 avdd.t93 dvss 2.10465f
C1870 avdd.n1038 dvss 1.34047f
C1871 avdd.n1040 dvss 0.196804f
C1872 avdd.n1041 dvss 0.196804f
C1873 avdd.t168 dvss 2.10465f
C1874 avdd.n1043 dvss 1.34047f
C1875 avdd.n1044 dvss 0.141631f
C1876 avdd.t144 dvss 2.10465f
C1877 avdd.n1046 dvss 1.34047f
C1878 avdd.n1047 dvss 0.141631f
C1879 avdd.n1048 dvss 0.141631f
C1880 avdd.n1049 dvss 1.34047f
C1881 avdd.n1051 dvss 0.196804f
C1882 avdd.t160 dvss 2.10465f
C1883 avdd.n1052 dvss 1.34047f
C1884 avdd.n1054 dvss 0.196804f
C1885 avdd.n1055 dvss 0.175474f
C1886 avdd.t109 dvss 2.10465f
C1887 avdd.n1057 dvss 1.34047f
C1888 avdd.n1058 dvss 0.120301f
C1889 avdd.n1059 dvss 0.257938f
C1890 avdd.n1060 dvss 0.927219f
C1891 avdd.n1061 dvss 0.900747f
C1892 avdd.n1062 dvss 0.179491f
C1893 avdd.n1063 dvss 0.206109f
C1894 avdd.n1064 dvss 0.78044f
C1895 avdd.n1065 dvss 0.301015f
C1896 avdd.n1066 dvss 0.140283f
C1897 avdd.n1067 dvss 0.259709f
C1898 avdd.t158 dvss 3.49651f
C1899 avdd.n1068 dvss 1.69278f
C1900 avdd.t159 dvss 0.120735f
C1901 avdd.n1070 dvss 0.968515f
C1902 avdd.n1071 dvss 1.97749f
C1903 avdd.n1072 dvss 2.43433f
C1904 avdd.n1073 dvss 1.94785f
C1905 avdd.n1074 dvss 1.05206f
C1906 avdd.n1075 dvss 1.07529f
C1907 avdd.n1076 dvss 4.644259f
C1908 avdd.n1077 dvss 4.644259f
C1909 avdd.n1078 dvss 17.7698f
C1910 avdd.n1079 dvss 4.61576f
C1911 avdd.n1080 dvss 17.3174f
C1912 avdd.n1081 dvss 17.7698f
C1913 avdd.n1082 dvss 17.3174f
C1914 avdd.n1083 dvss 4.61576f
C1915 avdd.n1084 dvss 1.08766f
C1916 avdd.n1085 dvss 1.08671f
C1917 avdd.n1086 dvss 1.07332f
C1918 avdd.n1087 dvss 0.257938f
C1919 avdd.n1089 dvss 0.175474f
C1920 avdd.n1091 dvss 0.196804f
C1921 avdd.n1093 dvss 0.196804f
C1922 avdd.n1095 dvss 0.196804f
C1923 avdd.n1097 dvss 0.196804f
C1924 avdd.n1099 dvss 0.196804f
C1925 avdd.n1101 dvss 0.196804f
C1926 avdd.n1103 dvss 0.196804f
C1927 avdd.n1105 dvss 0.195382f
C1928 avdd.t86 dvss 2.10465f
C1929 avdd.n1106 dvss 1.34047f
C1930 avdd.n1107 dvss 0.141631f
C1931 avdd.t113 dvss 2.10465f
C1932 avdd.n1108 dvss 1.34047f
C1933 avdd.n1109 dvss 0.141631f
C1934 avdd.t170 dvss 2.10465f
C1935 avdd.n1110 dvss 1.34047f
C1936 avdd.n1111 dvss 0.141631f
C1937 avdd.t95 dvss 2.10465f
C1938 avdd.n1112 dvss 1.34047f
C1939 avdd.n1113 dvss 0.141631f
C1940 avdd.t118 dvss 2.10465f
C1941 avdd.n1114 dvss 1.34047f
C1942 avdd.n1115 dvss 0.141631f
C1943 avdd.t146 dvss 2.10465f
C1944 avdd.n1116 dvss 1.34047f
C1945 avdd.n1117 dvss 0.141631f
C1946 avdd.t106 dvss 2.10465f
C1947 avdd.n1118 dvss 1.34047f
C1948 avdd.n1119 dvss 0.141631f
C1949 avdd.t128 dvss 2.10465f
C1950 avdd.n1120 dvss 1.34047f
C1951 avdd.n1121 dvss 0.140209f
C1952 avdd.t79 dvss 3.49651f
C1953 avdd.n1122 dvss 1.69278f
C1954 avdd.n1123 dvss 0.259709f
C1955 avdd.n1124 dvss 0.140283f
C1956 avdd.n1125 dvss 0.301015f
C1957 avdd.n1126 dvss 0.78044f
C1958 avdd.n1127 dvss 0.140283f
C1959 avdd.n1129 dvss 0.301791f
C1960 avdd.n1130 dvss 0.776758f
C1961 avdd.n1131 dvss 1.86745f
C1962 avdd.n1132 dvss 2.52205f
C1963 avdd.n1133 dvss 1.94784f
C1964 avdd.n1134 dvss 1.03703f
C1965 avdd.n1135 dvss 1.07017f
C1966 avdd.n1136 dvss 1.07332f
C1967 avdd.n1137 dvss 1.09835f
C1968 avdd.n1138 dvss 1.83172f
C1969 avdd.n1139 dvss 0.737267f
C1970 avdd.n1140 dvss 2.35767f
C1971 avdd.n1141 dvss 1.63565f
C1972 avdd.n1142 dvss 2.75705f
C1973 avdd.n1143 dvss 23.0904f
C1974 avdd.n1144 dvss 2.63303f
C1975 avdd.n1145 dvss 1.6959f
C1976 avdd.n1146 dvss 1.93486f
C1977 avdd.n1147 dvss 14.734401f
C1978 avdd.n1148 dvss 2.48436f
C1979 avdd.t340 dvss 1.62904f
C1980 avdd.t213 dvss 2.25453f
C1981 avdd.n1149 dvss 1.99568f
C1982 avdd.n1150 dvss 0.20375f
C1983 avdd.n1151 dvss 0.188858f
C1984 avdd.n1152 dvss 0.165742f
C1985 avdd.n1154 dvss 0.898386f
C1986 avdd.n1155 dvss 0.939824f
C1987 avdd.n1156 dvss 0.257938f
C1988 avdd.n1157 dvss 1.58216f
C1989 avdd.n1158 dvss 0.629059f
C1990 avdd.n1159 dvss 0.589894f
C1991 avdd.n1160 dvss 0.551818f
C1992 avdd.n1161 dvss 3.9961f
C1993 avdd.n1162 dvss 6.9044f
C1994 avdd.n1163 dvss 1.8298f
C1995 avdd.n1164 dvss 2.13126f
C1996 avdd.n1165 dvss 13.702299f
C1997 avdd.n1166 dvss 19.890001f
C1998 avdd.n1167 dvss 52.562603f
C1999 avdd.n1168 dvss 39.3676f
C2000 avdd.n1169 dvss 10.219099f
C2001 avdd.n1170 dvss 2.54131f
C2002 avdd.n1171 dvss 7.4696f
C2003 avdd.n1172 dvss 0.749362f
C2004 avdd.n1173 dvss 7.83749f
C2005 avdd.n1174 dvss 1.76577f
C2006 avdd.n1175 dvss 9.28326f
C2007 avdd.n1176 dvss 2.50544f
C2008 avdd.n1177 dvss 2.50732f
C2009 avdd.n1178 dvss 1.09589f
C2010 avdd.n1179 dvss 7.84177f
C2011 avdd.n1180 dvss 6.33529f
C2012 avdd.n1181 dvss 30.0285f
C2013 avdd.n1182 dvss 24.8949f
C2014 avdd.n1183 dvss 15.603301f
C2015 avdd.n1184 dvss 4.01126f
C2016 avdd.n1185 dvss 1.84112f
C2017 avdd.n1186 dvss 4.02745f
C2018 avdd.n1187 dvss 4.41765f
C2019 avdd.n1188 dvss 2.15978f
C2020 avdd.n1189 dvss 2.15723f
C2021 avdd.n1190 dvss 7.36437f
C2022 avdd.n1191 dvss 4.54554f
C2023 avdd.n1192 dvss 3.9387f
C2024 avdd.n1193 dvss 8.5683f
C2025 avdd.n1194 dvss 16.248499f
C2026 avdd.n1195 dvss 14.14f
C2027 avdd.n1196 dvss 6.48806f
C2028 avdd.n1197 dvss 14.127099f
C2029 avdd.n1198 dvss 54.3765f
C2030 avdd.n1199 dvss 76.4143f
C2031 avdd.n1200 dvss 75.227104f
C2032 avdd.n1201 dvss 19.551199f
C2033 avdd.n1202 dvss 1.58742f
C2034 avdd.n1203 dvss 1.94772f
C2035 avdd.n1204 dvss 1.79923f
C2036 avdd.n1205 dvss 3.99177f
C2037 avdd.n1206 dvss 33.806602f
C2038 avdd.n1207 dvss 55.4966f
C2039 avdd.n1208 dvss 2.37412f
C2040 avdd.t143 dvss 0.128868f
C2041 avdd.t202 dvss 0.128868f
C2042 avdd.n1209 dvss 0.327223f
C2043 avdd.n1210 dvss 0.730456f
C2044 avdd.n1211 dvss 1.81413f
C2045 avdd.n1212 dvss 1.695f
C2046 avdd.n1213 dvss 0.265705f
C2047 avdd.n1214 dvss 0.354515f
C2048 avdd.n1215 dvss 0.744085f
C2049 avdd.n1216 dvss 0.846264f
C2050 avdd.t425 dvss 5.64762f
C2051 avdd.t423 dvss 2.82381f
C2052 avdd.n1217 dvss 0.744085f
C2053 avdd.n1218 dvss 0.121474f
C2054 avdd.n1219 dvss 0.375451f
C2055 avdd.n1220 dvss 0.637382f
C2056 avdd.t426 dvss 6.20744f
C2057 avdd.t78 dvss 5.64762f
C2058 avdd.t428 dvss 5.64762f
C2059 avdd.t4 dvss 3.80739f
C2060 avdd.t421 dvss 3.5377f
C2061 avdd.n1221 dvss 0.346913f
C2062 avdd.n1222 dvss 8.3128f
C2063 avdd.t199 dvss 11.0573f
C2064 avdd.t122 dvss 7.265759f
C2065 avdd.t338 dvss 8.931499f
C2066 avdd.n1223 dvss 3.51487f
C2067 avdd.n1224 dvss 3.51487f
C2068 avdd.n1225 dvss 2.06209f
C2069 avdd.n1226 dvss 2.0377f
C2070 avdd.n1227 dvss 1.78233f
C2071 avdd.t203 dvss 4.31504f
C2072 avdd.t142 dvss 5.64762f
C2073 avdd.t201 dvss 5.64762f
C2074 avdd.t5 dvss 6.36151f
C2075 avdd.n1228 dvss 3.64875f
C2076 avdd.t48 dvss 8.10262f
C2077 avdd.t44 dvss 11.7863f
C2078 avdd.t46 dvss 12.155f
C2079 avdd.t50 dvss 9.11621f
C2080 avdd.n1229 dvss 6.07748f
C2081 avdd.t137 dvss 9.11621f
C2082 avdd.t362 dvss 12.155f
C2083 avdd.t364 dvss 12.155f
C2084 avdd.t154 dvss 12.155f
C2085 avdd.t366 dvss 12.155f
C2086 avdd.t368 dvss 12.155f
C2087 avdd.t99 dvss 10.2239f
C2088 avdd.n1230 dvss 8.71407f
C2089 avdd.n1231 dvss 1.05447f
C2090 avdd.n1232 dvss 1.06471f
C2091 avdd.n1233 dvss 3.59863f
C2092 avdd.t136 dvss 5.44629f
C2093 avdd.n1234 dvss 1.79091f
C2094 avdd.n1235 dvss 2.22604f
C2095 avdd.n1236 dvss 0.443709f
C2096 avdd.t101 dvss 0.477637f
C2097 avdd.t98 dvss 5.58077f
C2098 avdd.n1237 dvss 4.94641f
C2099 avdd.n1238 dvss 0.88709f
C2100 avdd.t369 dvss 0.128868f
C2101 avdd.t100 dvss 0.128868f
C2102 avdd.n1239 dvss 0.275381f
C2103 avdd.n1240 dvss 1.82615f
C2104 avdd.n1241 dvss 1.82615f
C2105 avdd.t365 dvss 0.128868f
C2106 avdd.t367 dvss 0.128868f
C2107 avdd.n1242 dvss 0.275381f
C2108 avdd.t155 dvss 0.257736f
C2109 avdd.n1243 dvss 0.265364f
C2110 avdd.t153 dvss 5.57075f
C2111 avdd.n1244 dvss 4.91093f
C2112 avdd.n1245 dvss 1.75079f
C2113 avdd.t51 dvss 0.128868f
C2114 avdd.n1246 dvss 0.262503f
C2115 avdd.t138 dvss 0.257736f
C2116 avdd.t363 dvss 0.128868f
C2117 avdd.n1247 dvss 0.275381f
C2118 avdd.n1248 dvss 1.8268f
C2119 avdd.n1249 dvss 1.25736f
C2120 avdd.n1250 dvss 0.208449f
C2121 avdd.n1251 dvss 2.21132f
C2122 avdd.n1252 dvss 1.76234f
C2123 avdd.n1253 dvss 1.75376f
C2124 avdd.t45 dvss 0.128868f
C2125 avdd.t47 dvss 0.128868f
C2126 avdd.n1254 dvss 0.275381f
C2127 avdd.n1255 dvss 1.7367f
C2128 avdd.t424 dvss 0.128868f
C2129 avdd.t49 dvss 0.128868f
C2130 avdd.n1256 dvss 0.275381f
C2131 avdd.n1257 dvss 2.39043f
C2132 avdd.n1258 dvss 1.82615f
C2133 avdd.t422 dvss 0.128868f
C2134 avdd.n1259 dvss 0.275381f
C2135 avdd.t123 dvss 0.606505f
C2136 avdd.t121 dvss 5.58077f
C2137 avdd.n1260 dvss 4.94641f
C2138 avdd.n1261 dvss 0.883188f
C2139 avdd.n1262 dvss 3.62799f
C2140 avdd.n1263 dvss 1.06471f
C2141 avdd.n1264 dvss 1.05447f
C2142 avdd.n1265 dvss 3.53886f
C2143 avdd.n1266 dvss 7.265759f
C2144 avdd.n1267 dvss 0.637382f
C2145 avdd.n1268 dvss 1.86976f
C2146 avdd.t205 dvss 0.539975f
C2147 avdd.n1269 dvss 1.33672f
C2148 avdd.t337 dvss 0.539975f
C2149 avdd.n1270 dvss 1.16514f
C2150 avdd.t141 dvss 1.07912f
C2151 avdd.n1271 dvss 0.978129f
C2152 avdd.t149 dvss 1.07897f
C2153 avdd.n1272 dvss 1.15815f
C2154 avdd.t77 dvss 1.07897f
C2155 avdd.n1273 dvss 1.30349f
C2156 avdd.n1274 dvss 0.199591f
C2157 avdd.n1275 dvss 0.604578f
C2158 avdd.t200 dvss 0.539975f
C2159 avdd.n1276 dvss 1.25984f
C2160 avdd.t335 dvss 0.128868f
C2161 avdd.t339 dvss 0.128868f
C2162 avdd.n1277 dvss 0.329341f
C2163 avdd.n1278 dvss 1.72572f
C2164 avdd.t347 dvss 0.128868f
C2165 avdd.t427 dvss 0.128868f
C2166 avdd.n1279 dvss 0.329341f
C2167 avdd.n1280 dvss 1.51264f
C2168 avdd.n1281 dvss 0.613128f
C2169 avdd.n1282 dvss 0.199591f
C2170 avdd.n1283 dvss 0.357819f
C2171 avdd.t131 dvss 1.74515f
C2172 avdd.n1284 dvss 3.63981f
C2173 avdd.t204 dvss 3.88785f
C2174 avdd.t346 dvss 5.81539f
C2175 avdd.n1285 dvss 0.121474f
C2176 avdd.n1286 dvss 0.346913f
C2177 avdd.n1287 dvss 4.43415f
C2178 avdd.t336 dvss 3.6904f
C2179 avdd.n1288 dvss 0.263845f
C2180 avdd.n1289 dvss 0.450444f
C2181 avdd.t132 dvss 3.65499f
C2182 avdd.n1290 dvss 0.450444f
C2183 avdd.n1291 dvss 0.809629f
C2184 avdd.n1292 dvss 0.345687f
C2185 avdd.n1293 dvss 0.19324f
C2186 avdd.n1294 dvss 0.25579f
C2187 avdd.n1295 dvss 0.659289f
C2188 avdd.t334 dvss 5.16112f
C2189 avdd.n1296 dvss 0.659289f
C2190 avdd.n1297 dvss 0.25579f
C2191 avdd.n1298 dvss 0.19324f
C2192 avdd.n1299 dvss 0.375451f
C2193 avdd.n1300 dvss 0.388199f
C2194 avdd.n1301 dvss 0.66168f
C2195 avdd.t150 dvss 4.1564f
C2196 avdd.n1302 dvss 0.66168f
C2197 avdd.n1303 dvss 0.366454f
C2198 avdd.n1304 dvss 0.285619f
C2199 avdd.n1305 dvss 1.86848f
C2200 avdd.n1306 dvss 2.71133f
C2201 avdd.n1307 dvss 18.0096f
C2202 avdd.n1308 dvss 37.8279f
C2203 avdd.n1309 dvss 24.6136f
C2204 avdd.t386 dvss 0.57241f
C2205 avdd.n1310 dvss 1.09164f
C2206 avdd.n1311 dvss 0.940945f
C2207 avdd.n1312 dvss 0.37963f
C2208 avdd.t400 dvss 0.128868f
C2209 avdd.t416 dvss 0.128868f
C2210 avdd.n1313 dvss 0.364688f
C2211 avdd.n1314 dvss 1.18763f
C2212 avdd.t396 dvss 0.128868f
C2213 avdd.t412 dvss 0.128868f
C2214 avdd.n1315 dvss 0.364688f
C2215 avdd.n1316 dvss 1.18763f
C2216 avdd.t408 dvss 0.128868f
C2217 avdd.t390 dvss 0.128868f
C2218 avdd.n1317 dvss 0.364688f
C2219 avdd.n1318 dvss 1.18763f
C2220 avdd.t404 dvss 0.128868f
C2221 avdd.t388 dvss 0.128868f
C2222 avdd.n1319 dvss 0.364688f
C2223 avdd.n1320 dvss 1.18763f
C2224 avdd.t402 dvss 0.128868f
C2225 avdd.t398 dvss 0.128868f
C2226 avdd.n1321 dvss 0.364688f
C2227 avdd.n1322 dvss 1.18763f
C2228 avdd.t414 dvss 0.128868f
C2229 avdd.t394 dvss 0.128868f
C2230 avdd.n1323 dvss 0.364688f
C2231 avdd.n1324 dvss 1.18763f
C2232 avdd.t410 dvss 0.128868f
C2233 avdd.t392 dvss 0.128868f
C2234 avdd.n1325 dvss 0.364688f
C2235 avdd.n1326 dvss 1.18763f
C2236 avdd.t406 dvss 0.57241f
C2237 avdd.n1327 dvss 1.26582f
C2238 avdd.n1328 dvss 1.24269f
C2239 avdd.n1329 dvss 0.389017f
C2240 avdd.n1330 dvss 1.14066f
C2241 avdd.n1331 dvss 0.37963f
C2242 avdd.n1332 dvss 0.550083f
C2243 avdd.n1333 dvss 1.14066f
C2244 avdd.n1334 dvss 3.74706f
C2245 avdd.t385 dvss 2.91873f
C2246 avdd.t399 dvss 2.41092f
C2247 avdd.t415 dvss 2.41092f
C2248 avdd.t395 dvss 2.41092f
C2249 avdd.t411 dvss 2.41092f
C2250 avdd.t407 dvss 2.41092f
C2251 avdd.t389 dvss 2.41092f
C2252 avdd.t403 dvss 1.80819f
C2253 avdd.n1335 dvss 1.20546f
C2254 avdd.t387 dvss 1.80819f
C2255 avdd.t401 dvss 2.41092f
C2256 avdd.t397 dvss 2.41092f
C2257 avdd.t413 dvss 2.41092f
C2258 avdd.t393 dvss 2.41092f
C2259 avdd.t409 dvss 2.41092f
C2260 avdd.t391 dvss 2.41092f
C2261 avdd.t405 dvss 2.91873f
C2262 avdd.n1336 dvss 3.74706f
C2263 avdd.n1337 dvss 0.389017f
C2264 avdd.n1338 dvss 0.670224f
C2265 avdd.n1339 dvss 1.32338f
C2266 avdd.n1340 dvss 1.24138f
C2267 avdd.n1341 dvss 0.451482f
C2268 avdd.n1342 dvss 1.68447f
C2269 avdd.n1343 dvss 1.42356f
C2270 avdd.n1344 dvss 1.33465f
C2271 avdd.n1345 dvss 2.21711f
C2272 avdd.n1346 dvss 1.33024f
C2273 avdd.n1347 dvss 0.775203f
C2274 avdd.n1348 dvss 0.193368f
C2275 avdd.n1349 dvss 5.17409f
C2276 avdd.t442 dvss 2.91873f
C2277 avdd.t441 dvss 2.41092f
C2278 avdd.t127 dvss 2.41092f
C2279 avdd.t434 dvss 2.41092f
C2280 avdd.t433 dvss 2.41092f
C2281 avdd.t90 dvss 2.41092f
C2282 avdd.t43 dvss 2.41092f
C2283 avdd.t42 dvss 2.41092f
C2284 avdd.t140 dvss 2.41092f
C2285 avdd.t212 dvss 2.41092f
C2286 avdd.t211 dvss 2.41092f
C2287 avdd.t112 dvss 2.41092f
C2288 avdd.t311 dvss 2.41092f
C2289 avdd.t312 dvss 2.41092f
C2290 avdd.t163 dvss 2.41092f
C2291 avdd.t323 dvss 2.41092f
C2292 avdd.t322 dvss 2.41092f
C2293 avdd.t103 dvss 2.41092f
C2294 avdd.t310 dvss 2.41092f
C2295 avdd.t309 dvss 2.41092f
C2296 avdd.t178 dvss 2.41092f
C2297 avdd.t349 dvss 2.41092f
C2298 avdd.t348 dvss 2.41092f
C2299 avdd.t167 dvss 2.41092f
C2300 avdd.t356 dvss 2.41092f
C2301 avdd.t357 dvss 2.41092f
C2302 avdd.t157 dvss 2.41092f
C2303 avdd.t436 dvss 2.41092f
C2304 avdd.t435 dvss 2.41092f
C2305 avdd.t165 dvss 2.41092f
C2306 avdd.t320 dvss 2.41092f
C2307 avdd.t321 dvss 2.41092f
C2308 avdd.t125 dvss 2.41092f
C2309 avdd.t439 dvss 2.41092f
C2310 avdd.t440 dvss 2.41092f
C2311 avdd.t176 dvss 2.41092f
C2312 avdd.t40 dvss 2.41092f
C2313 avdd.t41 dvss 2.41092f
C2314 avdd.t180 dvss 2.41092f
C2315 avdd.t375 dvss 2.41092f
C2316 avdd.t376 dvss 2.41092f
C2317 avdd.t152 dvss 2.41092f
C2318 avdd.t302 dvss 2.41092f
C2319 avdd.t301 dvss 2.41092f
C2320 avdd.t92 dvss 2.41092f
C2321 avdd.t262 dvss 2.41092f
C2322 avdd.t263 dvss 2.91873f
C2323 avdd.n1350 dvss 5.17409f
C2324 avdd.n1351 dvss 0.193725f
C2325 avdd.n1352 dvss 0.774242f
C2326 avdd.n1353 dvss 0.362835f
C2327 avdd.n1354 dvss 1.58506f
C2328 avdd.n1355 dvss 1.20551f
C2329 avss.t326 dvss 0.268751f
C2330 avss.n3 dvss 6.75695f
C2331 avss.n6 dvss 0.566482f
C2332 avss.n11 dvss 2.66222f
C2333 avss.t312 dvss 4.29356f
C2334 avss.t317 dvss 11.8082f
C2335 avss.n12 dvss 2.20901f
C2336 avss.n13 dvss 20.9681f
C2337 avss.n14 dvss 22.1122f
C2338 avss.n15 dvss 2.2117f
C2339 avss.n16 dvss 2.2104f
C2340 avss.n17 dvss 1.90754f
C2341 avss.n18 dvss 1.62554f
C2342 avss.n19 dvss 0.706789f
C2343 avss.n20 dvss 0.626109f
C2344 avss.t75 dvss 0.310265f
C2345 avss.n21 dvss 0.198678f
C2346 avss.n22 dvss 0.224592f
C2347 avss.n23 dvss 0.149121f
C2348 avss.n24 dvss 0.84204f
C2349 avss.n25 dvss 0.84204f
C2350 avss.t277 dvss 11.482599f
C2351 avss.t300 dvss 11.8082f
C2352 avss.t154 dvss 11.8082f
C2353 avss.t337 dvss 11.8082f
C2354 avss.t376 dvss 11.8082f
C2355 avss.t306 dvss 11.8082f
C2356 avss.t237 dvss 11.8082f
C2357 avss.t296 dvss 11.8082f
C2358 avss.t271 dvss 11.8082f
C2359 avss.t242 dvss 11.8082f
C2360 avss.t262 dvss 11.8082f
C2361 avss.t261 dvss 11.8082f
C2362 avss.t270 dvss 11.8082f
C2363 avss.t216 dvss 11.8082f
C2364 avss.t382 dvss 11.8082f
C2365 avss.t257 dvss 11.8082f
C2366 avss.t354 dvss 11.8082f
C2367 avss.t318 dvss 11.8082f
C2368 avss.t4 dvss 5.94733f
C2369 avss.n26 dvss 13.411599f
C2370 avss.n44 dvss 0.332218f
C2371 avss.n45 dvss 0.326909f
C2372 avss.n60 dvss 0.332218f
C2373 avss.n61 dvss 0.326909f
C2374 avss.n76 dvss 0.332218f
C2375 avss.n77 dvss 0.326909f
C2376 avss.n92 dvss 0.332218f
C2377 avss.n93 dvss 0.326909f
C2378 avss.n108 dvss 0.332218f
C2379 avss.n109 dvss 0.326909f
C2380 avss.n124 dvss 0.332218f
C2381 avss.n125 dvss 0.326909f
C2382 avss.n140 dvss 0.332218f
C2383 avss.n141 dvss 0.326909f
C2384 avss.n149 dvss 0.401577f
C2385 avss.n153 dvss 0.419945f
C2386 avss.n161 dvss 0.326909f
C2387 avss.n162 dvss 0.332218f
C2388 avss.n175 dvss 0.326909f
C2389 avss.n176 dvss 0.332218f
C2390 avss.n189 dvss 0.326909f
C2391 avss.n190 dvss 0.332218f
C2392 avss.n203 dvss 0.326909f
C2393 avss.n204 dvss 0.332218f
C2394 avss.n217 dvss 0.326909f
C2395 avss.n218 dvss 0.332218f
C2396 avss.n231 dvss 0.326909f
C2397 avss.n232 dvss 0.332218f
C2398 avss.n245 dvss 0.326909f
C2399 avss.n246 dvss 0.332218f
C2400 avss.n259 dvss 0.326909f
C2401 avss.n260 dvss 0.332218f
C2402 avss.n266 dvss 0.799724f
C2403 avss.n267 dvss 20.7399f
C2404 avss.t328 dvss 6.15926f
C2405 avss.t297 dvss 6.15926f
C2406 avss.t152 dvss 6.15926f
C2407 avss.t55 dvss 6.15926f
C2408 avss.t331 dvss 6.15926f
C2409 avss.t258 dvss 6.15926f
C2410 avss.t56 dvss 6.15926f
C2411 avss.t19 dvss 6.56811f
C2412 avss.n268 dvss 3.91016f
C2413 avss.t298 dvss 3.45257f
C2414 avss.n269 dvss 0.250887f
C2415 avss.n270 dvss 0.186167f
C2416 avss.n271 dvss 0.1132f
C2417 avss.n272 dvss 0.131097f
C2418 avss.n273 dvss 0.215339f
C2419 avss.n274 dvss 1.41349f
C2420 avss.n275 dvss 1.26024f
C2421 avss.n276 dvss 1.07892f
C2422 avss.t80 dvss 0.310248f
C2423 avss.t135 dvss 0.310248f
C2424 avss.t129 dvss 0.310265f
C2425 avss.n277 dvss 0.1925f
C2426 avss.n278 dvss 0.185709f
C2427 avss.t122 dvss 0.310265f
C2428 avss.n279 dvss 0.19255f
C2429 avss.t131 dvss 0.310265f
C2430 avss.n280 dvss 0.190331f
C2431 avss.t127 dvss 0.310265f
C2432 avss.n281 dvss 0.190464f
C2433 avss.t104 dvss 0.310265f
C2434 avss.n282 dvss 0.190702f
C2435 avss.t84 dvss 0.310265f
C2436 avss.n283 dvss 0.154735f
C2437 avss.t63 dvss 0.310265f
C2438 avss.n285 dvss 0.189612f
C2439 avss.n286 dvss 0.18568f
C2440 avss.t86 dvss 0.310265f
C2441 avss.n287 dvss 0.19255f
C2442 avss.t67 dvss 0.310265f
C2443 avss.n288 dvss 0.190331f
C2444 avss.t115 dvss 0.310265f
C2445 avss.n289 dvss 0.190331f
C2446 avss.t82 dvss 0.310265f
C2447 avss.n290 dvss 0.190331f
C2448 avss.t108 dvss 0.310265f
C2449 avss.n291 dvss 0.199473f
C2450 avss.n292 dvss 0.641703f
C2451 avss.n293 dvss 9.78569f
C2452 avss.n294 dvss 0.773733f
C2453 avss.n295 dvss 1.02802f
C2454 avss.t110 dvss 4.09377f
C2455 avss.t112 dvss 0.158938f
C2456 avss.n296 dvss 1.54547f
C2457 avss.n297 dvss 0.401096f
C2458 avss.n298 dvss 0.197936f
C2459 avss.n299 dvss 0.163183f
C2460 avss.n300 dvss 1.25443f
C2461 avss.n301 dvss 1.25443f
C2462 avss.t88 dvss 4.09377f
C2463 avss.n302 dvss 0.163183f
C2464 avss.t89 dvss 0.201402f
C2465 avss.n303 dvss 1.54547f
C2466 avss.n304 dvss 0.45849f
C2467 avss.n305 dvss 0.502647f
C2468 avss.n306 dvss 0.692104f
C2469 avss.n307 dvss 0.692104f
C2470 avss.n308 dvss 1.09153f
C2471 avss.n309 dvss 1.09153f
C2472 avss.t213 dvss 4.40637f
C2473 avss.t320 dvss 3.69892f
C2474 avss.n310 dvss 0.451633f
C2475 avss.n311 dvss 0.22261f
C2476 avss.n312 dvss 0.45849f
C2477 avss.t93 dvss 4.09377f
C2478 avss.n313 dvss 1.54547f
C2479 avss.t94 dvss 0.201402f
C2480 avss.n314 dvss 0.163183f
C2481 avss.n315 dvss 1.25443f
C2482 avss.n316 dvss 0.163183f
C2483 avss.n317 dvss 1.25443f
C2484 avss.t71 dvss 4.09377f
C2485 avss.t74 dvss 0.158938f
C2486 avss.n318 dvss 1.54547f
C2487 avss.n319 dvss 0.401096f
C2488 avss.n320 dvss 2.02822f
C2489 avss.t65 dvss 0.349415f
C2490 avss.n321 dvss 0.64704f
C2491 avss.n322 dvss 0.128891f
C2492 avss.n323 dvss 0.149988f
C2493 avss.n324 dvss 0.399555f
C2494 avss.n325 dvss 0.399555f
C2495 avss.t163 dvss 4.91169f
C2496 avss.t295 dvss 3.59786f
C2497 avss.t107 dvss 5.8819f
C2498 avss.t164 dvss 5.35636f
C2499 avss.t299 dvss 3.59786f
C2500 avss.t134 dvss 4.10318f
C2501 avss.t285 dvss 3.59786f
C2502 avss.t360 dvss 3.53722f
C2503 avss.t5 dvss 3.59786f
C2504 avss.t66 dvss 4.99254f
C2505 avss.t174 dvss 6.24572f
C2506 avss.t18 dvss 3.59786f
C2507 avss.t243 dvss 5.13402f
C2508 avss.n326 dvss 0.78405f
C2509 avss.n327 dvss 0.78405f
C2510 avss.n328 dvss 0.405117f
C2511 avss.n329 dvss 0.836963f
C2512 avss.n330 dvss 0.676102f
C2513 avss.n331 dvss 0.588602f
C2514 avss.n332 dvss 0.783978f
C2515 avss.n333 dvss 0.798746f
C2516 avss.n334 dvss 0.702705f
C2517 avss.t92 dvss 0.154277f
C2518 avss.t90 dvss 1.81398f
C2519 avss.n335 dvss 1.6064f
C2520 avss.n336 dvss 0.707168f
C2521 avss.n337 dvss 0.627132f
C2522 avss.n338 dvss 0.662218f
C2523 avss.n339 dvss 0.367097f
C2524 avss.n340 dvss 0.38026f
C2525 avss.n341 dvss 0.647338f
C2526 avss.n342 dvss 0.647338f
C2527 avss.t69 dvss 2.32303f
C2528 avss.n343 dvss 1.85321f
C2529 avss.t121 dvss 0.154277f
C2530 avss.t119 dvss 1.81398f
C2531 avss.n344 dvss 1.6064f
C2532 avss.n345 dvss 0.705217f
C2533 avss.n346 dvss 0.351612f
C2534 avss.n347 dvss 0.682669f
C2535 avss.n348 dvss 0.203433f
C2536 avss.n349 dvss 0.19684f
C2537 avss.n350 dvss 17.9279f
C2538 avss.t120 dvss 4.55932f
C2539 avss.t44 dvss 4.96505f
C2540 avss.t45 dvss 4.62363f
C2541 avss.t218 dvss 7.6404f
C2542 avss.t380 dvss 7.6404f
C2543 avss.t17 dvss 7.6404f
C2544 avss.t314 dvss 7.6404f
C2545 avss.t206 dvss 7.6404f
C2546 avss.t308 dvss 7.6404f
C2547 avss.t339 dvss 7.6404f
C2548 avss.t263 dvss 7.6404f
C2549 avss.t253 dvss 7.6404f
C2550 avss.t377 dvss 7.6404f
C2551 avss.t204 dvss 7.6404f
C2552 avss.t24 dvss 7.6404f
C2553 avss.t315 dvss 7.6404f
C2554 avss.t275 dvss 7.6404f
C2555 avss.t199 dvss 7.6404f
C2556 avss.t338 dvss 7.6404f
C2557 avss.t329 dvss 3.37552f
C2558 avss.t20 dvss 14.9866f
C2559 avss.t230 dvss 15.2808f
C2560 avss.t341 dvss 7.66061f
C2561 avss.n351 dvss 5.154241f
C2562 avss.t355 dvss 7.62019f
C2563 avss.t273 dvss 7.6404f
C2564 avss.t309 dvss 7.6404f
C2565 avss.t205 dvss 7.6404f
C2566 avss.t59 dvss 7.6404f
C2567 avss.t280 dvss 7.6404f
C2568 avss.t15 dvss 7.6404f
C2569 avss.t245 dvss 7.6404f
C2570 avss.t319 dvss 7.6404f
C2571 avss.t370 dvss 7.6404f
C2572 avss.t305 dvss 7.6404f
C2573 avss.t47 dvss 7.6404f
C2574 avss.t352 dvss 7.6404f
C2575 avss.t334 dvss 7.6404f
C2576 avss.t252 dvss 7.6404f
C2577 avss.t178 dvss 7.6404f
C2578 avss.t177 dvss 7.6404f
C2579 avss.t219 dvss 7.6404f
C2580 avss.t381 dvss 7.6404f
C2581 avss.t301 dvss 3.8202f
C2582 avss.n352 dvss 5.154241f
C2583 avss.t307 dvss 6.30636f
C2584 avss.t54 dvss 6.75104f
C2585 avss.n353 dvss 7.63676f
C2586 avss.t70 dvss 1.51324f
C2587 avss.n354 dvss 2.48252f
C2588 avss.t25 dvss 3.79323f
C2589 avss.t43 dvss 4.96505f
C2590 avss.t91 dvss 4.1115f
C2591 avss.n355 dvss 32.3852f
C2592 avss.t181 dvss 0.795915f
C2593 avss.n356 dvss 0.207329f
C2594 avss.n357 dvss 0.207329f
C2595 avss.t96 dvss 7.05778f
C2596 avss.n360 dvss 0.938161f
C2597 avss.n361 dvss 0.938161f
C2598 avss.n363 dvss 0.296614f
C2599 avss.n364 dvss 0.57227f
C2600 avss.n365 dvss 0.469902f
C2601 avss.n366 dvss 0.469902f
C2602 avss.n367 dvss 2.15938f
C2603 avss.n368 dvss 0.468647f
C2604 avss.n369 dvss 0.262958f
C2605 avss.n370 dvss 1.2431f
C2606 avss.n373 dvss 0.203226f
C2607 avss.n377 dvss 0.203754f
C2608 avss.n379 dvss 0.111489f
C2609 avss.n381 dvss 0.113557f
C2610 avss.n382 dvss 0.109193f
C2611 avss.n383 dvss 0.129041f
C2612 avss.n384 dvss 0.514356f
C2613 avss.n385 dvss 1.0014f
C2614 avss.t26 dvss 0.65894f
C2615 avss.t28 dvss 0.377405f
C2616 avss.t32 dvss 0.377405f
C2617 avss.t38 dvss 0.377405f
C2618 avss.t30 dvss 0.283051f
C2619 avss.n386 dvss 0.47633f
C2620 avss.n387 dvss 0.58503f
C2621 avss.n388 dvss 0.349486f
C2622 avss.n389 dvss 0.392198f
C2623 avss.n390 dvss 0.78405f
C2624 avss.n391 dvss 0.78405f
C2625 avss.t378 dvss 11.8082f
C2626 avss.t357 dvss 11.8082f
C2627 avss.t58 dvss 11.8082f
C2628 avss.t23 dvss 11.673f
C2629 avss.t336 dvss 14.0232f
C2630 avss.t316 dvss 5.31594f
C2631 avss.n392 dvss 0.206798f
C2632 avss.n393 dvss 0.206798f
C2633 avss.n394 dvss 0.29074f
C2634 avss.t137 dvss 0.456853f
C2635 avss.t159 dvss 1.65744f
C2636 avss.n395 dvss 5.21488f
C2637 avss.t138 dvss 5.98296f
C2638 avss.t353 dvss 5.21488f
C2639 avss.t324 dvss 7.6404f
C2640 avss.t379 dvss 5.31594f
C2641 avss.t198 dvss 7.33721f
C2642 avss.n396 dvss 0.294947f
C2643 avss.n397 dvss 0.294947f
C2644 avss.n398 dvss 0.173184f
C2645 avss.n399 dvss 0.144197f
C2646 avss.t160 dvss 0.217588f
C2647 avss.t325 dvss 0.213102f
C2648 avss.n400 dvss 0.868457f
C2649 avss.t133 dvss 0.349431f
C2650 avss.n401 dvss 0.296889f
C2651 avss.t106 dvss 0.349412f
C2652 avss.n402 dvss 0.342553f
C2653 avss.n403 dvss 0.205284f
C2654 avss.t161 dvss 7.6404f
C2655 avss.t310 dvss 9.25742f
C2656 avss.t2 dvss 7.6404f
C2657 avss.t57 dvss 4.62871f
C2658 avss.n404 dvss 7.6404f
C2659 avss.t231 dvss 4.62871f
C2660 avss.t0 dvss 7.6404f
C2661 avss.t259 dvss 7.62019f
C2662 avss.t283 dvss 2.78935f
C2663 avss.t358 dvss 6.488279f
C2664 avss.t346 dvss 7.33721f
C2665 avss.n405 dvss 5.154241f
C2666 avss.n406 dvss 5.86168f
C2667 avss.n407 dvss 0.297166f
C2668 avss.n409 dvss 0.120103f
C2669 avss.n410 dvss 0.109931f
C2670 avss.t359 dvss 0.213102f
C2671 avss.n411 dvss 0.418376f
C2672 avss.n412 dvss 0.156149f
C2673 avss.n413 dvss 0.560087f
C2674 avss.t162 dvss 0.213102f
C2675 avss.n414 dvss 0.418593f
C2676 avss.n415 dvss 0.155007f
C2677 avss.n416 dvss 0.120103f
C2678 avss.n418 dvss 0.297166f
C2679 avss.n419 dvss 1.79893f
C2680 avss.t61 dvss 4.87126f
C2681 avss.n420 dvss 5.84147f
C2682 avss.n421 dvss 0.205609f
C2683 avss.n422 dvss 0.113389f
C2684 avss.n423 dvss 0.299297f
C2685 avss.n424 dvss 0.113887f
C2686 avss.n425 dvss 0.205609f
C2687 avss.n426 dvss 7.6404f
C2688 avss.t185 dvss 10.5106f
C2689 avss.t311 dvss 8.61061f
C2690 avss.n427 dvss 25.4096f
C2691 avss.n428 dvss 0.273716f
C2692 avss.n429 dvss 0.39203f
C2693 avss.n430 dvss 0.897599f
C2694 avss.n431 dvss 1.08082f
C2695 avss.n432 dvss 0.95396f
C2696 avss.n433 dvss 0.705031f
C2697 avss.n434 dvss 0.781633f
C2698 avss.n435 dvss 27.925001f
C2699 avss.t274 dvss 10.2316f
C2700 avss.t335 dvss 10.808599f
C2701 avss.t361 dvss 10.808599f
C2702 avss.t153 dvss 10.808599f
C2703 avss.t304 dvss 10.808599f
C2704 avss.t330 dvss 10.808599f
C2705 avss.t21 dvss 9.00716f
C2706 avss.n436 dvss 15.096701f
C2707 avss.t42 dvss 7.20572f
C2708 avss.t332 dvss 10.808599f
C2709 avss.t214 dvss 8.10644f
C2710 avss.n437 dvss 5.40429f
C2711 avss.t345 dvss 8.10644f
C2712 avss.t46 dvss 10.808599f
C2713 avss.t254 dvss 10.808599f
C2714 avss.t303 dvss 10.808599f
C2715 avss.t251 dvss 10.808599f
C2716 avss.t281 dvss 10.808599f
C2717 avss.t272 dvss 10.808599f
C2718 avss.t207 dvss 10.808599f
C2719 avss.t220 dvss 10.808599f
C2720 avss.t6 dvss 9.03575f
C2721 avss.n438 dvss 8.921371f
C2722 avss.n439 dvss 0.783978f
C2723 avss.n440 dvss 0.118969f
C2724 avss.n441 dvss 0.134237f
C2725 avss.n442 dvss 0.307129f
C2726 avss.n443 dvss 0.27886f
C2727 avss.n444 dvss 0.104223f
C2728 avss.n446 dvss 0.215561f
C2729 avss.t211 dvss 0.955458f
C2730 avss.t188 dvss 8.929259f
C2731 avss.t190 dvss 6.69694f
C2732 avss.n448 dvss 4.46463f
C2733 avss.t192 dvss 6.69694f
C2734 avss.t186 dvss 8.929259f
C2735 avss.t78 dvss 7.05778f
C2736 avss.n449 dvss 0.946545f
C2737 avss.n450 dvss 2.97088f
C2738 avss.n451 dvss 0.244143f
C2739 avss.t209 dvss 0.286975f
C2740 avss.t40 dvss 0.377405f
C2741 avss.t36 dvss 0.377405f
C2742 avss.t34 dvss 0.283051f
C2743 avss.n452 dvss 0.110247f
C2744 avss.n453 dvss 0.215561f
C2745 avss.n455 dvss 0.104223f
C2746 avss.n456 dvss 0.191958f
C2747 avss.n457 dvss 1.16186f
C2748 avss.t99 dvss 1.11622f
C2749 avss.t77 dvss 1.11622f
C2750 avss.n458 dvss 0.552993f
C2751 avss.n460 dvss 0.135342f
C2752 avss.n461 dvss 0.124977f
C2753 avss.n463 dvss 0.552993f
C2754 avss.n466 dvss 0.262958f
C2755 avss.n467 dvss 0.262958f
C2756 avss.n468 dvss 0.138191f
C2757 avss.t399 dvss 0.739019f
C2758 avss.n469 dvss 0.508077f
C2759 avss.t400 dvss 0.739019f
C2760 avss.n470 dvss 0.314947f
C2761 avss.t397 dvss 0.739019f
C2762 avss.n471 dvss 0.314947f
C2763 avss.t398 dvss 0.739019f
C2764 avss.n472 dvss 0.314947f
C2765 avss.t396 dvss 0.739019f
C2766 avss.n473 dvss 0.314947f
C2767 avss.t391 dvss 0.739019f
C2768 avss.n474 dvss 0.314947f
C2769 avss.t392 dvss 0.739019f
C2770 avss.n475 dvss 0.314947f
C2771 avss.t388 dvss 0.739019f
C2772 avss.n476 dvss 1.27942f
C2773 avss.t113 dvss 0.703139f
C2774 avss.n507 dvss 0.320366f
C2775 avss.n508 dvss 0.565285f
C2776 avss.n509 dvss 0.130132f
C2777 avss.n510 dvss 0.565934f
C2778 avss.n511 dvss 0.130035f
C2779 avss.n512 dvss 0.565934f
C2780 avss.n513 dvss 0.565934f
C2781 avss.n514 dvss 2.06477f
C2782 avss.n515 dvss 0.130332f
C2783 avss.n516 dvss 0.260088f
C2784 avss.n517 dvss 0.566164f
C2785 avss.n518 dvss 2.07947f
C2786 avss.n519 dvss 2.06477f
C2787 avss.n520 dvss 2.07947f
C2788 avss.n521 dvss 0.566164f
C2789 avss.n522 dvss 0.259687f
C2790 avss.n523 dvss 0.130033f
C2791 avss.n524 dvss 0.528695f
C2792 avss.n525 dvss 0.364911f
C2793 avss.n530 dvss 0.174247f
C2794 avss.n532 dvss 0.227005f
C2795 avss.t114 dvss 1.16359f
C2796 avss.n538 dvss 0.725466f
C2797 avss.n544 dvss 0.17126f
C2798 avss.n548 dvss 1.55227f
C2799 avss.n552 dvss 0.174247f
C2800 avss.n555 dvss 0.237026f
C2801 avss.n557 dvss 0.237026f
C2802 avss.n563 dvss 0.174247f
C2803 avss.n564 dvss 0.780568f
C2804 avss.n571 dvss 0.232964f
C2805 avss.n572 dvss 0.232964f
C2806 avss.n573 dvss 0.17126f
C2807 avss.n580 dvss 0.749429f
C2808 avss.n581 dvss 0.22294f
C2809 avss.n582 dvss 1.4441f
C2810 avss.n588 dvss 0.22294f
C2811 avss.n589 dvss 1.41775f
C2812 avss.n597 dvss 0.166879f
C2813 avss.n598 dvss 0.166879f
C2814 avss.n599 dvss 0.227005f
C2815 avss.n605 dvss 1.49876f
C2816 avss.n606 dvss 0.771646f
C2817 avss.n607 dvss 0.174247f
C2818 avss.n611 dvss 0.119914f
C2819 avss.n612 dvss 3.59244f
C2820 avss.n613 dvss 0.20945f
C2821 avss.n614 dvss 0.100509f
C2822 avss.n615 dvss 0.111514f
C2823 avss.n616 dvss 0.310785f
C2824 avss.n617 dvss 11.381599f
C2825 avss.n618 dvss 13.5304f
C2826 avss.n619 dvss 3.86195f
C2827 avss.t385 dvss 0.734641f
C2828 avss.n620 dvss 0.372042f
C2829 avss.t387 dvss 0.734641f
C2830 avss.n621 dvss 0.309894f
C2831 avss.t386 dvss 0.734641f
C2832 avss.n622 dvss 0.309894f
C2833 avss.t389 dvss 0.734641f
C2834 avss.n623 dvss 0.309894f
C2835 avss.t393 dvss 0.734641f
C2836 avss.n624 dvss 0.309894f
C2837 avss.t390 dvss 0.734641f
C2838 avss.n625 dvss 0.309894f
C2839 avss.t395 dvss 0.734641f
C2840 avss.n626 dvss 0.309894f
C2841 avss.t394 dvss 0.734641f
C2842 avss.n627 dvss 0.506256f
C2843 avss.n628 dvss 0.14152f
C2844 avss.t95 dvss 1.11622f
C2845 avss.n629 dvss 0.552993f
C2846 avss.t124 dvss 1.11622f
C2847 avss.n631 dvss 0.552993f
C2848 avss.n634 dvss 0.262958f
C2849 avss.n636 dvss 0.135342f
C2850 avss.n638 dvss 0.124977f
C2851 avss.n639 dvss 0.468647f
C2852 avss.n640 dvss 0.538393f
C2853 avss.n641 dvss 0.621504f
C2854 avss.n646 dvss 0.135342f
C2855 avss.n647 dvss 0.625278f
C2856 avss.n648 dvss 0.538394f
C2857 avss.n649 dvss 0.296614f
C2858 avss.n651 dvss 0.946545f
C2859 avss.n652 dvss 2.84896f
C2860 avss.n653 dvss 1.37135f
C2861 avss.t183 dvss 2.159f
C2862 avss.t179 dvss 1.21267f
C2863 avss.n654 dvss 1.11553f
C2864 avss.t321 dvss 2.13393f
C2865 avss.t323 dvss 2.03366f
C2866 avss.n655 dvss 27.431501f
C2867 avss.n656 dvss 0.212891f
C2868 avss.n657 dvss 0.124131f
C2869 avss.n658 dvss 0.122205f
C2870 avss.n660 dvss 0.212891f
C2871 avss.n661 dvss 12.0911f
C2872 avss.n662 dvss 45.845398f
C2873 avss.n663 dvss 15.4238f
C2874 avss.n664 dvss 0.653748f
C2875 avss.n665 dvss 0.19684f
C2876 avss.n666 dvss 0.203433f
C2877 avss.n667 dvss 0.682669f
C2878 avss.n668 dvss 0.494072f
C2879 avss.t356 dvss 0.233402f
C2880 avss.n669 dvss 1.07607f
C2881 avss.n670 dvss 0.713059f
C2882 avss.n671 dvss 0.963873f
C2883 avss.n672 dvss 0.704934f
C2884 avss.n673 dvss 0.789014f
C2885 avss.n674 dvss 0.582393f
C2886 avss.n675 dvss 0.405117f
C2887 avss.n676 dvss 0.393574f
C2888 avss.n677 dvss 0.783978f
C2889 avss.n678 dvss 7.6404f
C2890 avss.t282 dvss 12.6329f
C2891 avss.t208 dvss 11.6829f
C2892 avss.n679 dvss 7.6404f
C2893 avss.t236 dvss 7.55955f
C2894 avss.n680 dvss 7.6404f
C2895 avss.t147 dvss 4.507431f
C2896 avss.t172 dvss 4.42658f
C2897 avss.t169 dvss 6.81168f
C2898 avss.t176 dvss 3.59786f
C2899 avss.t175 dvss 0.586168f
C2900 avss.t72 dvss 3.59786f
C2901 avss.t166 dvss 6.99359f
C2902 avss.t167 dvss 3.6585f
C2903 avss.t225 dvss 3.59786f
C2904 avss.t168 dvss 7.13508f
C2905 avss.t170 dvss 4.10318f
C2906 avss.t215 dvss 3.59786f
C2907 avss.t171 dvss 6.6904f
C2908 avss.n681 dvss 0.128891f
C2909 avss.n682 dvss 0.232286f
C2910 avss.n683 dvss 0.395365f
C2911 avss.t173 dvss 4.54786f
C2912 avss.n684 dvss 0.395365f
C2913 avss.n685 dvss 0.203313f
C2914 avss.n686 dvss 0.149988f
C2915 avss.n687 dvss 0.859294f
C2916 avss.n688 dvss 1.08621f
C2917 avss.n689 dvss 1.02802f
C2918 avss.n690 dvss 0.271068f
C2919 avss.t101 dvss 4.09377f
C2920 avss.t103 dvss 0.158938f
C2921 avss.n691 dvss 1.54547f
C2922 avss.n692 dvss 0.401096f
C2923 avss.n693 dvss 0.163183f
C2924 avss.n694 dvss 1.25443f
C2925 avss.n695 dvss 1.25443f
C2926 avss.t117 dvss 4.09377f
C2927 avss.n696 dvss 0.163183f
C2928 avss.t118 dvss 0.201402f
C2929 avss.n697 dvss 1.54547f
C2930 avss.n698 dvss 0.45849f
C2931 avss.n699 dvss 0.198368f
C2932 avss.n702 dvss 0.150988f
C2933 avss.n703 dvss 0.271068f
C2934 avss.t142 dvss 4.09377f
C2935 avss.t144 dvss 0.158938f
C2936 avss.n704 dvss 1.54547f
C2937 avss.n705 dvss 0.401096f
C2938 avss.n706 dvss 0.163183f
C2939 avss.n707 dvss 1.25443f
C2940 avss.n708 dvss 1.25443f
C2941 avss.t60 dvss 4.09377f
C2942 avss.n709 dvss 0.163183f
C2943 avss.t62 dvss 0.201402f
C2944 avss.n710 dvss 1.54547f
C2945 avss.n711 dvss 0.45849f
C2946 avss.n712 dvss 0.151419f
C2947 avss.n713 dvss 0.223041f
C2948 avss.n714 dvss 0.45849f
C2949 avss.t145 dvss 4.09377f
C2950 avss.n715 dvss 1.54547f
C2951 avss.t146 dvss 0.201402f
C2952 avss.n716 dvss 0.163183f
C2953 avss.n717 dvss 1.25443f
C2954 avss.n718 dvss 0.163183f
C2955 avss.n719 dvss 1.25443f
C2956 avss.t139 dvss 4.09377f
C2957 avss.t141 dvss 0.158938f
C2958 avss.n720 dvss 1.54547f
C2959 avss.n721 dvss 0.401096f
C2960 avss.n722 dvss 0.271068f
C2961 avss.n723 dvss 1.02802f
C2962 avss.n724 dvss 1.04748f
C2963 avss.n725 dvss 0.271068f
C2964 avss.n726 dvss 0.451201f
C2965 avss.n727 dvss 0.640078f
C2966 avss.n728 dvss 0.644263f
C2967 avss.n729 dvss 1.09076f
C2968 avss.n730 dvss 2.72871f
C2969 avss.n731 dvss 1.09076f
C2970 avss.n732 dvss 0.642533f
C2971 avss.n733 dvss 0.744592f
C2972 avss.n734 dvss 0.502216f
C2973 avss.n735 dvss 0.271068f
C2974 avss.n736 dvss 0.923217f
C2975 avss.n737 dvss 0.731243f
C2976 avss.n738 dvss 7.71343f
C2977 avss.n739 dvss 4.79285f
C2978 avss.n740 dvss 0.131959f
C2979 avss.n741 dvss 0.608012f
C2980 avss.n742 dvss 0.144664f
C2981 avss.n743 dvss 0.28472f
C2982 avss.n744 dvss 0.849372f
C2983 avss.n745 dvss 3.86116f
C2984 avss.t244 dvss 2.27788f
C2985 avss.t349 dvss 3.65686f
C2986 avss.t350 dvss 2.02251f
C2987 avss.t276 dvss 1.81822f
C2988 avss.t109 dvss 3.43214f
C2989 avss.t371 dvss 2.24723f
C2990 avss.t260 dvss 1.81822f
C2991 avss.t372 dvss 3.20742f
C2992 avss.t83 dvss 2.47196f
C2993 avss.t302 dvss 1.81822f
C2994 avss.t238 dvss 2.98269f
C2995 avss.t239 dvss 2.69668f
C2996 avss.t313 dvss 1.81822f
C2997 avss.t116 dvss 2.75797f
C2998 avss.t10 dvss 2.92141f
C2999 avss.t383 dvss 1.81822f
C3000 avss.t7 dvss 2.53325f
C3001 avss.t68 dvss 3.14613f
C3002 avss.t375 dvss 1.81822f
C3003 avss.t49 dvss 2.30852f
C3004 avss.t50 dvss 3.37085f
C3005 avss.t16 dvss 1.81822f
C3006 avss.t87 dvss 2.0838f
C3007 avss.t203 dvss 3.59558f
C3008 avss.t340 dvss 1.81822f
C3009 avss.t200 dvss 1.85908f
C3010 avss.t81 dvss 3.63643f
C3011 avss.t196 dvss 2.00208f
C3012 avss.t351 dvss 1.81822f
C3013 avss.t197 dvss 3.45257f
C3014 avss.t64 dvss 2.22681f
C3015 avss.t255 dvss 1.81822f
C3016 avss.t269 dvss 3.22785f
C3017 avss.t266 dvss 2.45153f
C3018 avss.t279 dvss 1.81822f
C3019 avss.t85 dvss 3.00312f
C3020 avss.t156 dvss 2.67625f
C3021 avss.t246 dvss 1.81822f
C3022 avss.t155 dvss 2.7784f
C3023 avss.t105 dvss 2.90098f
C3024 avss.t384 dvss 1.81822f
C3025 avss.t224 dvss 2.55368f
C3026 avss.t221 dvss 3.1257f
C3027 avss.t22 dvss 1.81822f
C3028 avss.t128 dvss 2.32895f
C3029 avss.t14 dvss 3.35042f
C3030 avss.t217 dvss 1.81822f
C3031 avss.t13 dvss 2.10423f
C3032 avss.t132 dvss 3.57515f
C3033 avss.t264 dvss 1.81822f
C3034 avss.t366 dvss 1.87951f
C3035 avss.t369 dvss 3.63643f
C3036 avss.t123 dvss 1.98165f
C3037 avss.t53 dvss 1.81822f
C3038 avss.t235 dvss 3.473f
C3039 avss.t232 dvss 2.20638f
C3040 avss.t165 dvss 1.81822f
C3041 avss.t136 dvss 3.24828f
C3042 avss.t364 dvss 2.4311f
C3043 avss.t256 dvss 1.81822f
C3044 avss.t365 dvss 3.02355f
C3045 avss.t130 dvss 2.65582f
C3046 avss.t344 dvss 1.81822f
C3047 avss.t226 dvss 2.79883f
C3048 avss.t227 dvss 2.88055f
C3049 avss.t265 dvss 1.81822f
C3050 avss.t76 dvss 2.57411f
C3051 avss.t149 dvss 3.10527f
C3052 avss.t333 dvss 1.81822f
C3053 avss.t148 dvss 2.80904f
C3054 avss.n746 dvss 3.24828f
C3055 avss.n747 dvss 0.849372f
C3056 avss.n749 dvss 0.256662f
C3057 avss.n751 dvss 1.08758f
C3058 avss.n752 dvss 2.76626f
C3059 avss.t278 dvss 0.227476f
C3060 avss.n753 dvss 3.91401f
C3061 avss.n754 dvss 1.82249f
C3062 avss.n755 dvss 2.20901f
C3063 avss.n756 dvss 3.48781f
C3064 avss.n757 dvss 3.64219f
C3065 avss.n758 dvss 2.16255f
C3066 avss.n759 dvss 1.1045f
C3067 avss.n760 dvss 1.1058f
C3068 avss.n761 dvss 2.20901f
C3069 avss.t48 dvss 9.48092f
C3070 avss.n762 dvss 15.612599f
C3071 avss.n763 dvss 12.200099f
C3072 avss.t342 dvss 2.75655f
C3073 avss.n769 dvss 0.157327f
C3074 avss.n770 dvss 0.330781f
C3075 avss.n775 dvss 0.213402f
C3076 rstring_mux_0.vtrip12.n2 dvss 0.516678f
C3077 rstring_mux_0.vtrip12.n3 dvss 1.03041f
C3078 rstring_mux_0.vtrip12.t2 dvss 0.287839f
C3079 vin.n0 dvss 0.390096f
C3080 vin.n1 dvss 0.182832f
C3081 vin.n2 dvss 0.179545f
C3082 vin.t30 dvss 0.137532f
C3083 vin.n3 dvss 0.16178f
C3084 vin.n4 dvss 0.440394f
C3085 vin.n5 dvss 0.379768f
C3086 vin.n6 dvss 0.179545f
C3087 vin.t71 dvss 0.137532f
C3088 vin.n7 dvss 0.16178f
C3089 vin.n8 dvss 0.440394f
C3090 vin.n9 dvss 0.440394f
C3091 vin.n10 dvss 0.440394f
C3092 vin.n11 dvss 0.440394f
C3093 vin.n12 dvss 0.440394f
C3094 vin.n13 dvss 0.440394f
C3095 vin.n14 dvss 0.440394f
C3096 vin.n15 dvss 0.440394f
C3097 vin.n16 dvss 0.440394f
C3098 vin.n17 dvss 0.440394f
C3099 vin.n18 dvss 0.440394f
C3100 vin.n19 dvss 0.440394f
C3101 vin.t20 dvss 0.291564f
C3102 vin.n20 dvss 0.405281f
C3103 vin.n21 dvss 0.16178f
C3104 vin.t76 dvss 0.137532f
C3105 vin.n22 dvss 0.179545f
C3106 vin.n23 dvss 0.379768f
C3107 vin.n24 dvss 0.182832f
C3108 vin.n25 dvss 0.16178f
C3109 vin.t74 dvss 0.137532f
C3110 vin.n26 dvss 0.179545f
C3111 vin.n27 dvss 0.379768f
C3112 vin.n28 dvss 0.182832f
C3113 vin.n29 dvss 0.16178f
C3114 vin.t32 dvss 0.137532f
C3115 vin.n30 dvss 0.179545f
C3116 vin.n31 dvss 0.379768f
C3117 vin.n32 dvss 0.182832f
C3118 vin.n33 dvss 0.16178f
C3119 vin.t41 dvss 0.137532f
C3120 vin.n34 dvss 0.179545f
C3121 vin.n35 dvss 0.379768f
C3122 vin.n36 dvss 0.182832f
C3123 vin.n37 dvss 0.16178f
C3124 vin.t39 dvss 0.137532f
C3125 vin.n38 dvss 0.179545f
C3126 vin.n39 dvss 0.379768f
C3127 vin.n40 dvss 0.182832f
C3128 vin.n41 dvss 0.16178f
C3129 vin.t73 dvss 0.137532f
C3130 vin.n42 dvss 0.179545f
C3131 vin.n43 dvss 0.379768f
C3132 vin.n44 dvss 0.182832f
C3133 vin.n45 dvss 0.16178f
C3134 vin.t75 dvss 0.137532f
C3135 vin.n46 dvss 0.179545f
C3136 vin.n47 dvss 0.379768f
C3137 vin.n48 dvss 0.182832f
C3138 vin.n49 dvss 0.16178f
C3139 vin.t77 dvss 0.137532f
C3140 vin.n50 dvss 0.179545f
C3141 vin.n51 dvss 0.379768f
C3142 vin.n52 dvss 0.182832f
C3143 vin.n53 dvss 0.16178f
C3144 vin.t40 dvss 0.137532f
C3145 vin.n54 dvss 0.179545f
C3146 vin.n55 dvss 0.379768f
C3147 vin.n56 dvss 0.182832f
C3148 vin.n57 dvss 0.16178f
C3149 vin.t42 dvss 0.137532f
C3150 vin.n58 dvss 0.179545f
C3151 vin.n59 dvss 0.379768f
C3152 vin.n60 dvss 0.182832f
C3153 vin.n61 dvss 0.16178f
C3154 vin.t72 dvss 0.137532f
C3155 vin.n62 dvss 0.179545f
C3156 vin.n63 dvss 0.379768f
C3157 vin.n64 dvss 0.182832f
C3158 vin.t101 dvss 1.11409f
C3159 vin.t104 dvss 1.01142f
C3160 vin.n65 dvss 1.32508f
C3161 vin.t103 dvss 1.11409f
C3162 vin.t108 dvss 1.01142f
C3163 vin.n66 dvss 1.32062f
C3164 vin.t102 dvss 1.11409f
C3165 vin.t107 dvss 1.01142f
C3166 vin.n68 dvss 1.32062f
C3167 vin.t105 dvss 1.11409f
C3168 vin.t96 dvss 1.01142f
C3169 vin.n70 dvss 1.32062f
C3170 vin.t109 dvss 1.11409f
C3171 vin.t98 dvss 1.01142f
C3172 vin.n72 dvss 1.32062f
C3173 vin.t106 dvss 1.11409f
C3174 vin.t97 dvss 1.01142f
C3175 vin.n74 dvss 1.32062f
C3176 vin.t95 dvss 1.11409f
C3177 vin.t100 dvss 1.01142f
C3178 vin.n76 dvss 1.32062f
C3179 vin.t94 dvss 1.11409f
C3180 vin.t99 dvss 1.01142f
C3181 vin.n78 dvss 1.32062f
C3182 vin.n79 dvss 3.52016f
C3183 vin.n80 dvss 5.25466f
C3184 vin.n81 dvss 0.182832f
C3185 vin.n82 dvss 0.379768f
C3186 vin.n83 dvss 0.179545f
C3187 vin.t31 dvss 0.137532f
C3188 vin.n84 dvss 0.16178f
C3189 vin.n85 dvss 0.440394f
C3190 vin.t69 dvss 0.312823f
C3191 vin.n86 dvss 0.843292f
C3192 vin.n87 dvss 0.204863f
C3193 vin.t34 dvss 0.137532f
C3194 vin.n88 dvss 0.220707f
C3195 vin.n89 dvss 0.797877f
C3196 vin.n90 dvss 0.204863f
C3197 vin.t66 dvss 0.137532f
C3198 vin.n91 dvss 0.220707f
C3199 vin.n92 dvss 0.797877f
C3200 vin.n93 dvss 0.204863f
C3201 vin.t35 dvss 0.137532f
C3202 vin.n94 dvss 0.220707f
C3203 vin.n95 dvss 0.797877f
C3204 vin.n96 dvss 0.204863f
C3205 vin.t63 dvss 0.137532f
C3206 vin.n97 dvss 0.220707f
C3207 vin.n98 dvss 0.797877f
C3208 vin.n99 dvss 0.204863f
C3209 vin.t68 dvss 0.137532f
C3210 vin.n100 dvss 0.220707f
C3211 vin.n101 dvss 0.797877f
C3212 vin.n102 dvss 0.204863f
C3213 vin.t65 dvss 0.137532f
C3214 vin.n103 dvss 0.220707f
C3215 vin.n104 dvss 0.797877f
C3216 vin.n105 dvss 0.204863f
C3217 vin.t93 dvss 0.137532f
C3218 vin.n106 dvss 0.220707f
C3219 vin.n107 dvss 0.797877f
C3220 vin.n108 dvss 0.204863f
C3221 vin.t67 dvss 0.137532f
C3222 vin.n109 dvss 0.220707f
C3223 vin.n110 dvss 0.797877f
C3224 vin.n111 dvss 0.204863f
C3225 vin.t33 dvss 0.137532f
C3226 vin.n112 dvss 0.220707f
C3227 vin.n113 dvss 0.797877f
C3228 vin.n114 dvss 0.204863f
C3229 vin.t43 dvss 0.137532f
C3230 vin.n115 dvss 0.220707f
C3231 vin.n116 dvss 0.797877f
C3232 vin.n117 dvss 0.204863f
C3233 vin.t45 dvss 0.137532f
C3234 vin.n118 dvss 0.220707f
C3235 vin.n119 dvss 0.797877f
C3236 vin.n120 dvss 0.204863f
C3237 vin.t36 dvss 0.137532f
C3238 vin.n121 dvss 0.220707f
C3239 vin.n122 dvss 0.797877f
C3240 vin.n123 dvss 0.204863f
C3241 vin.t46 dvss 0.137532f
C3242 vin.n124 dvss 0.220707f
C3243 vin.n125 dvss 0.797877f
C3244 vin.n126 dvss 0.204863f
C3245 vin.t44 dvss 0.137532f
C3246 vin.n127 dvss 0.220707f
C3247 vin.t92 dvss 0.274286f
C3248 vin.n128 dvss 0.46542f
C3249 vin.t10 dvss 0.297788f
C3250 vin.n129 dvss 0.842484f
C3251 vin.n130 dvss 0.220707f
C3252 vin.t64 dvss 0.137532f
C3253 vin.n131 dvss 0.204863f
C3254 vin.n132 dvss 0.797877f
C3255 vin.n133 dvss 0.179545f
C3256 vin.t78 dvss 0.137532f
C3257 vin.n134 dvss 0.16178f
C3258 vin.n135 dvss 0.440394f
C3259 vin.n136 dvss 0.379768f
C3260 vin.n137 dvss 0.11545f
.ends

