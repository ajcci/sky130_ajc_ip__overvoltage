magic
tech sky130A
magscale 1 2
timestamp 1712077413
<< nwell >>
rect -3232 -797 3232 797
<< mvpmos >>
rect -2974 -500 -2174 500
rect -2116 -500 -1316 500
rect -1258 -500 -458 500
rect -400 -500 400 500
rect 458 -500 1258 500
rect 1316 -500 2116 500
rect 2174 -500 2974 500
<< mvpdiff >>
rect -3032 488 -2974 500
rect -3032 -488 -3020 488
rect -2986 -488 -2974 488
rect -3032 -500 -2974 -488
rect -2174 488 -2116 500
rect -2174 -488 -2162 488
rect -2128 -488 -2116 488
rect -2174 -500 -2116 -488
rect -1316 488 -1258 500
rect -1316 -488 -1304 488
rect -1270 -488 -1258 488
rect -1316 -500 -1258 -488
rect -458 488 -400 500
rect -458 -488 -446 488
rect -412 -488 -400 488
rect -458 -500 -400 -488
rect 400 488 458 500
rect 400 -488 412 488
rect 446 -488 458 488
rect 400 -500 458 -488
rect 1258 488 1316 500
rect 1258 -488 1270 488
rect 1304 -488 1316 488
rect 1258 -500 1316 -488
rect 2116 488 2174 500
rect 2116 -488 2128 488
rect 2162 -488 2174 488
rect 2116 -500 2174 -488
rect 2974 488 3032 500
rect 2974 -488 2986 488
rect 3020 -488 3032 488
rect 2974 -500 3032 -488
<< mvpdiffc >>
rect -3020 -488 -2986 488
rect -2162 -488 -2128 488
rect -1304 -488 -1270 488
rect -446 -488 -412 488
rect 412 -488 446 488
rect 1270 -488 1304 488
rect 2128 -488 2162 488
rect 2986 -488 3020 488
<< mvnsubdiff >>
rect -3166 719 3166 731
rect -3166 685 -3058 719
rect 3058 685 3166 719
rect -3166 673 3166 685
rect -3166 623 -3108 673
rect -3166 -623 -3154 623
rect -3120 -623 -3108 623
rect 3108 623 3166 673
rect -3166 -673 -3108 -623
rect 3108 -623 3120 623
rect 3154 -623 3166 623
rect 3108 -673 3166 -623
rect -3166 -685 3166 -673
rect -3166 -719 -3058 -685
rect 3058 -719 3166 -685
rect -3166 -731 3166 -719
<< mvnsubdiffcont >>
rect -3058 685 3058 719
rect -3154 -623 -3120 623
rect 3120 -623 3154 623
rect -3058 -719 3058 -685
<< poly >>
rect -2974 581 -2174 597
rect -2974 547 -2958 581
rect -2190 547 -2174 581
rect -2974 500 -2174 547
rect -2116 581 -1316 597
rect -2116 547 -2100 581
rect -1332 547 -1316 581
rect -2116 500 -1316 547
rect -1258 581 -458 597
rect -1258 547 -1242 581
rect -474 547 -458 581
rect -1258 500 -458 547
rect -400 581 400 597
rect -400 547 -384 581
rect 384 547 400 581
rect -400 500 400 547
rect 458 581 1258 597
rect 458 547 474 581
rect 1242 547 1258 581
rect 458 500 1258 547
rect 1316 581 2116 597
rect 1316 547 1332 581
rect 2100 547 2116 581
rect 1316 500 2116 547
rect 2174 581 2974 597
rect 2174 547 2190 581
rect 2958 547 2974 581
rect 2174 500 2974 547
rect -2974 -547 -2174 -500
rect -2974 -581 -2958 -547
rect -2190 -581 -2174 -547
rect -2974 -597 -2174 -581
rect -2116 -547 -1316 -500
rect -2116 -581 -2100 -547
rect -1332 -581 -1316 -547
rect -2116 -597 -1316 -581
rect -1258 -547 -458 -500
rect -1258 -581 -1242 -547
rect -474 -581 -458 -547
rect -1258 -597 -458 -581
rect -400 -547 400 -500
rect -400 -581 -384 -547
rect 384 -581 400 -547
rect -400 -597 400 -581
rect 458 -547 1258 -500
rect 458 -581 474 -547
rect 1242 -581 1258 -547
rect 458 -597 1258 -581
rect 1316 -547 2116 -500
rect 1316 -581 1332 -547
rect 2100 -581 2116 -547
rect 1316 -597 2116 -581
rect 2174 -547 2974 -500
rect 2174 -581 2190 -547
rect 2958 -581 2974 -547
rect 2174 -597 2974 -581
<< polycont >>
rect -2958 547 -2190 581
rect -2100 547 -1332 581
rect -1242 547 -474 581
rect -384 547 384 581
rect 474 547 1242 581
rect 1332 547 2100 581
rect 2190 547 2958 581
rect -2958 -581 -2190 -547
rect -2100 -581 -1332 -547
rect -1242 -581 -474 -547
rect -384 -581 384 -547
rect 474 -581 1242 -547
rect 1332 -581 2100 -547
rect 2190 -581 2958 -547
<< locali >>
rect -3154 685 -3058 719
rect 3058 685 3154 719
rect -3154 623 -3120 685
rect 3120 623 3154 685
rect -2974 547 -2958 581
rect -2190 547 -2174 581
rect -2116 547 -2100 581
rect -1332 547 -1316 581
rect -1258 547 -1242 581
rect -474 547 -458 581
rect -400 547 -384 581
rect 384 547 400 581
rect 458 547 474 581
rect 1242 547 1258 581
rect 1316 547 1332 581
rect 2100 547 2116 581
rect 2174 547 2190 581
rect 2958 547 2974 581
rect -3020 488 -2986 504
rect -3020 -504 -2986 -488
rect -2162 488 -2128 504
rect -2162 -504 -2128 -488
rect -1304 488 -1270 504
rect -1304 -504 -1270 -488
rect -446 488 -412 504
rect -446 -504 -412 -488
rect 412 488 446 504
rect 412 -504 446 -488
rect 1270 488 1304 504
rect 1270 -504 1304 -488
rect 2128 488 2162 504
rect 2128 -504 2162 -488
rect 2986 488 3020 504
rect 2986 -504 3020 -488
rect -2974 -581 -2958 -547
rect -2190 -581 -2174 -547
rect -2116 -581 -2100 -547
rect -1332 -581 -1316 -547
rect -1258 -581 -1242 -547
rect -474 -581 -458 -547
rect -400 -581 -384 -547
rect 384 -581 400 -547
rect 458 -581 474 -547
rect 1242 -581 1258 -547
rect 1316 -581 1332 -547
rect 2100 -581 2116 -547
rect 2174 -581 2190 -547
rect 2958 -581 2974 -547
rect -3154 -685 -3120 -623
rect 3120 -685 3154 -623
rect -3154 -719 -3058 -685
rect 3058 -719 3154 -685
<< viali >>
rect -2958 547 -2190 581
rect -2100 547 -1332 581
rect -1242 547 -474 581
rect -384 547 384 581
rect 474 547 1242 581
rect 1332 547 2100 581
rect 2190 547 2958 581
rect -3020 -488 -2986 488
rect -2162 -488 -2128 488
rect -1304 -488 -1270 488
rect -446 -488 -412 488
rect 412 -488 446 488
rect 1270 -488 1304 488
rect 2128 -488 2162 488
rect 2986 -488 3020 488
rect -2958 -581 -2190 -547
rect -2100 -581 -1332 -547
rect -1242 -581 -474 -547
rect -384 -581 384 -547
rect 474 -581 1242 -547
rect 1332 -581 2100 -547
rect 2190 -581 2958 -547
<< metal1 >>
rect -2970 581 -2178 587
rect -2970 547 -2958 581
rect -2190 547 -2178 581
rect -2970 541 -2178 547
rect -2112 581 -1320 587
rect -2112 547 -2100 581
rect -1332 547 -1320 581
rect -2112 541 -1320 547
rect -1254 581 -462 587
rect -1254 547 -1242 581
rect -474 547 -462 581
rect -1254 541 -462 547
rect -396 581 396 587
rect -396 547 -384 581
rect 384 547 396 581
rect -396 541 396 547
rect 462 581 1254 587
rect 462 547 474 581
rect 1242 547 1254 581
rect 462 541 1254 547
rect 1320 581 2112 587
rect 1320 547 1332 581
rect 2100 547 2112 581
rect 1320 541 2112 547
rect 2178 581 2970 587
rect 2178 547 2190 581
rect 2958 547 2970 581
rect 2178 541 2970 547
rect -3026 488 -2980 500
rect -3026 -488 -3020 488
rect -2986 -488 -2980 488
rect -3026 -500 -2980 -488
rect -2168 488 -2122 500
rect -2168 -488 -2162 488
rect -2128 -488 -2122 488
rect -2168 -500 -2122 -488
rect -1310 488 -1264 500
rect -1310 -488 -1304 488
rect -1270 -488 -1264 488
rect -1310 -500 -1264 -488
rect -452 488 -406 500
rect -452 -488 -446 488
rect -412 -488 -406 488
rect -452 -500 -406 -488
rect 406 488 452 500
rect 406 -488 412 488
rect 446 -488 452 488
rect 406 -500 452 -488
rect 1264 488 1310 500
rect 1264 -488 1270 488
rect 1304 -488 1310 488
rect 1264 -500 1310 -488
rect 2122 488 2168 500
rect 2122 -488 2128 488
rect 2162 -488 2168 488
rect 2122 -500 2168 -488
rect 2980 488 3026 500
rect 2980 -488 2986 488
rect 3020 -488 3026 488
rect 2980 -500 3026 -488
rect -2970 -547 -2178 -541
rect -2970 -581 -2958 -547
rect -2190 -581 -2178 -547
rect -2970 -587 -2178 -581
rect -2112 -547 -1320 -541
rect -2112 -581 -2100 -547
rect -1332 -581 -1320 -547
rect -2112 -587 -1320 -581
rect -1254 -547 -462 -541
rect -1254 -581 -1242 -547
rect -474 -581 -462 -547
rect -1254 -587 -462 -581
rect -396 -547 396 -541
rect -396 -581 -384 -547
rect 384 -581 396 -547
rect -396 -587 396 -581
rect 462 -547 1254 -541
rect 462 -581 474 -547
rect 1242 -581 1254 -547
rect 462 -587 1254 -581
rect 1320 -547 2112 -541
rect 1320 -581 1332 -547
rect 2100 -581 2112 -547
rect 1320 -587 2112 -581
rect 2178 -547 2970 -541
rect 2178 -581 2190 -547
rect 2958 -581 2970 -547
rect 2178 -587 2970 -581
<< properties >>
string FIXED_BBOX -3137 -702 3137 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 4 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
