magic
tech sky130A
magscale 1 2
timestamp 1712109191
<< nwell >>
rect -1030 -797 1030 797
<< mvpmos >>
rect -772 -500 -652 500
rect -594 -500 -474 500
rect -416 -500 -296 500
rect -238 -500 -118 500
rect -60 -500 60 500
rect 118 -500 238 500
rect 296 -500 416 500
rect 474 -500 594 500
rect 652 -500 772 500
<< mvpdiff >>
rect -830 488 -772 500
rect -830 -488 -818 488
rect -784 -488 -772 488
rect -830 -500 -772 -488
rect -652 488 -594 500
rect -652 -488 -640 488
rect -606 -488 -594 488
rect -652 -500 -594 -488
rect -474 488 -416 500
rect -474 -488 -462 488
rect -428 -488 -416 488
rect -474 -500 -416 -488
rect -296 488 -238 500
rect -296 -488 -284 488
rect -250 -488 -238 488
rect -296 -500 -238 -488
rect -118 488 -60 500
rect -118 -488 -106 488
rect -72 -488 -60 488
rect -118 -500 -60 -488
rect 60 488 118 500
rect 60 -488 72 488
rect 106 -488 118 488
rect 60 -500 118 -488
rect 238 488 296 500
rect 238 -488 250 488
rect 284 -488 296 488
rect 238 -500 296 -488
rect 416 488 474 500
rect 416 -488 428 488
rect 462 -488 474 488
rect 416 -500 474 -488
rect 594 488 652 500
rect 594 -488 606 488
rect 640 -488 652 488
rect 594 -500 652 -488
rect 772 488 830 500
rect 772 -488 784 488
rect 818 -488 830 488
rect 772 -500 830 -488
<< mvpdiffc >>
rect -818 -488 -784 488
rect -640 -488 -606 488
rect -462 -488 -428 488
rect -284 -488 -250 488
rect -106 -488 -72 488
rect 72 -488 106 488
rect 250 -488 284 488
rect 428 -488 462 488
rect 606 -488 640 488
rect 784 -488 818 488
<< mvnsubdiff >>
rect -964 719 964 731
rect -964 685 -856 719
rect 856 685 964 719
rect -964 673 964 685
rect -964 623 -906 673
rect -964 -623 -952 623
rect -918 -623 -906 623
rect 906 623 964 673
rect -964 -673 -906 -623
rect 906 -623 918 623
rect 952 -623 964 623
rect 906 -673 964 -623
rect -964 -685 964 -673
rect -964 -719 -856 -685
rect 856 -719 964 -685
rect -964 -731 964 -719
<< mvnsubdiffcont >>
rect -856 685 856 719
rect -952 -623 -918 623
rect 918 -623 952 623
rect -856 -719 856 -685
<< poly >>
rect -772 581 -652 597
rect -772 547 -756 581
rect -668 547 -652 581
rect -772 500 -652 547
rect -594 581 -474 597
rect -594 547 -578 581
rect -490 547 -474 581
rect -594 500 -474 547
rect -416 581 -296 597
rect -416 547 -400 581
rect -312 547 -296 581
rect -416 500 -296 547
rect -238 581 -118 597
rect -238 547 -222 581
rect -134 547 -118 581
rect -238 500 -118 547
rect -60 581 60 597
rect -60 547 -44 581
rect 44 547 60 581
rect -60 500 60 547
rect 118 581 238 597
rect 118 547 134 581
rect 222 547 238 581
rect 118 500 238 547
rect 296 581 416 597
rect 296 547 312 581
rect 400 547 416 581
rect 296 500 416 547
rect 474 581 594 597
rect 474 547 490 581
rect 578 547 594 581
rect 474 500 594 547
rect 652 581 772 597
rect 652 547 668 581
rect 756 547 772 581
rect 652 500 772 547
rect -772 -547 -652 -500
rect -772 -581 -756 -547
rect -668 -581 -652 -547
rect -772 -597 -652 -581
rect -594 -547 -474 -500
rect -594 -581 -578 -547
rect -490 -581 -474 -547
rect -594 -597 -474 -581
rect -416 -547 -296 -500
rect -416 -581 -400 -547
rect -312 -581 -296 -547
rect -416 -597 -296 -581
rect -238 -547 -118 -500
rect -238 -581 -222 -547
rect -134 -581 -118 -547
rect -238 -597 -118 -581
rect -60 -547 60 -500
rect -60 -581 -44 -547
rect 44 -581 60 -547
rect -60 -597 60 -581
rect 118 -547 238 -500
rect 118 -581 134 -547
rect 222 -581 238 -547
rect 118 -597 238 -581
rect 296 -547 416 -500
rect 296 -581 312 -547
rect 400 -581 416 -547
rect 296 -597 416 -581
rect 474 -547 594 -500
rect 474 -581 490 -547
rect 578 -581 594 -547
rect 474 -597 594 -581
rect 652 -547 772 -500
rect 652 -581 668 -547
rect 756 -581 772 -547
rect 652 -597 772 -581
<< polycont >>
rect -756 547 -668 581
rect -578 547 -490 581
rect -400 547 -312 581
rect -222 547 -134 581
rect -44 547 44 581
rect 134 547 222 581
rect 312 547 400 581
rect 490 547 578 581
rect 668 547 756 581
rect -756 -581 -668 -547
rect -578 -581 -490 -547
rect -400 -581 -312 -547
rect -222 -581 -134 -547
rect -44 -581 44 -547
rect 134 -581 222 -547
rect 312 -581 400 -547
rect 490 -581 578 -547
rect 668 -581 756 -547
<< locali >>
rect -952 685 -856 719
rect 856 685 952 719
rect -952 623 -918 685
rect 918 623 952 685
rect -772 547 -756 581
rect -668 547 -652 581
rect -594 547 -578 581
rect -490 547 -474 581
rect -416 547 -400 581
rect -312 547 -296 581
rect -238 547 -222 581
rect -134 547 -118 581
rect -60 547 -44 581
rect 44 547 60 581
rect 118 547 134 581
rect 222 547 238 581
rect 296 547 312 581
rect 400 547 416 581
rect 474 547 490 581
rect 578 547 594 581
rect 652 547 668 581
rect 756 547 772 581
rect -818 488 -784 504
rect -818 -504 -784 -488
rect -640 488 -606 504
rect -640 -504 -606 -488
rect -462 488 -428 504
rect -462 -504 -428 -488
rect -284 488 -250 504
rect -284 -504 -250 -488
rect -106 488 -72 504
rect -106 -504 -72 -488
rect 72 488 106 504
rect 72 -504 106 -488
rect 250 488 284 504
rect 250 -504 284 -488
rect 428 488 462 504
rect 428 -504 462 -488
rect 606 488 640 504
rect 606 -504 640 -488
rect 784 488 818 504
rect 784 -504 818 -488
rect -772 -581 -756 -547
rect -668 -581 -652 -547
rect -594 -581 -578 -547
rect -490 -581 -474 -547
rect -416 -581 -400 -547
rect -312 -581 -296 -547
rect -238 -581 -222 -547
rect -134 -581 -118 -547
rect -60 -581 -44 -547
rect 44 -581 60 -547
rect 118 -581 134 -547
rect 222 -581 238 -547
rect 296 -581 312 -547
rect 400 -581 416 -547
rect 474 -581 490 -547
rect 578 -581 594 -547
rect 652 -581 668 -547
rect 756 -581 772 -547
rect -952 -685 -918 -623
rect 918 -685 952 -623
rect -952 -719 -856 -685
rect 856 -719 952 -685
<< viali >>
rect -756 547 -668 581
rect -578 547 -490 581
rect -400 547 -312 581
rect -222 547 -134 581
rect -44 547 44 581
rect 134 547 222 581
rect 312 547 400 581
rect 490 547 578 581
rect 668 547 756 581
rect -818 -488 -784 488
rect -640 -488 -606 488
rect -462 -488 -428 488
rect -284 -488 -250 488
rect -106 -488 -72 488
rect 72 -488 106 488
rect 250 -488 284 488
rect 428 -488 462 488
rect 606 -488 640 488
rect 784 -488 818 488
rect -756 -581 -668 -547
rect -578 -581 -490 -547
rect -400 -581 -312 -547
rect -222 -581 -134 -547
rect -44 -581 44 -547
rect 134 -581 222 -547
rect 312 -581 400 -547
rect 490 -581 578 -547
rect 668 -581 756 -547
<< metal1 >>
rect -768 581 -656 587
rect -768 547 -756 581
rect -668 547 -656 581
rect -768 541 -656 547
rect -590 581 -478 587
rect -590 547 -578 581
rect -490 547 -478 581
rect -590 541 -478 547
rect -412 581 -300 587
rect -412 547 -400 581
rect -312 547 -300 581
rect -412 541 -300 547
rect -234 581 -122 587
rect -234 547 -222 581
rect -134 547 -122 581
rect -234 541 -122 547
rect -56 581 56 587
rect -56 547 -44 581
rect 44 547 56 581
rect -56 541 56 547
rect 122 581 234 587
rect 122 547 134 581
rect 222 547 234 581
rect 122 541 234 547
rect 300 581 412 587
rect 300 547 312 581
rect 400 547 412 581
rect 300 541 412 547
rect 478 581 590 587
rect 478 547 490 581
rect 578 547 590 581
rect 478 541 590 547
rect 656 581 768 587
rect 656 547 668 581
rect 756 547 768 581
rect 656 541 768 547
rect -824 488 -778 500
rect -824 -488 -818 488
rect -784 -488 -778 488
rect -824 -500 -778 -488
rect -646 488 -600 500
rect -646 -488 -640 488
rect -606 -488 -600 488
rect -646 -500 -600 -488
rect -468 488 -422 500
rect -468 -488 -462 488
rect -428 -488 -422 488
rect -468 -500 -422 -488
rect -290 488 -244 500
rect -290 -488 -284 488
rect -250 -488 -244 488
rect -290 -500 -244 -488
rect -112 488 -66 500
rect -112 -488 -106 488
rect -72 -488 -66 488
rect -112 -500 -66 -488
rect 66 488 112 500
rect 66 -488 72 488
rect 106 -488 112 488
rect 66 -500 112 -488
rect 244 488 290 500
rect 244 -488 250 488
rect 284 -488 290 488
rect 244 -500 290 -488
rect 422 488 468 500
rect 422 -488 428 488
rect 462 -488 468 488
rect 422 -500 468 -488
rect 600 488 646 500
rect 600 -488 606 488
rect 640 -488 646 488
rect 600 -500 646 -488
rect 778 488 824 500
rect 778 -488 784 488
rect 818 -488 824 488
rect 778 -500 824 -488
rect -768 -547 -656 -541
rect -768 -581 -756 -547
rect -668 -581 -656 -547
rect -768 -587 -656 -581
rect -590 -547 -478 -541
rect -590 -581 -578 -547
rect -490 -581 -478 -547
rect -590 -587 -478 -581
rect -412 -547 -300 -541
rect -412 -581 -400 -547
rect -312 -581 -300 -547
rect -412 -587 -300 -581
rect -234 -547 -122 -541
rect -234 -581 -222 -547
rect -134 -581 -122 -547
rect -234 -587 -122 -581
rect -56 -547 56 -541
rect -56 -581 -44 -547
rect 44 -581 56 -547
rect -56 -587 56 -581
rect 122 -547 234 -541
rect 122 -581 134 -547
rect 222 -581 234 -547
rect 122 -587 234 -581
rect 300 -547 412 -541
rect 300 -581 312 -547
rect 400 -581 412 -547
rect 300 -587 412 -581
rect 478 -547 590 -541
rect 478 -581 490 -547
rect 578 -581 590 -547
rect 478 -587 590 -581
rect 656 -547 768 -541
rect 656 -581 668 -547
rect 756 -581 768 -547
rect 656 -587 768 -581
<< properties >>
string FIXED_BBOX -935 -702 935 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.6 m 1 nf 9 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
