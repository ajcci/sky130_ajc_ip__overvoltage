magic
tech sky130A
magscale 1 2
timestamp 1712339160
<< error_p >>
rect -4444 1342 -4370 1351
rect -4444 1286 -4435 1342
rect -4444 1277 -4370 1286
rect -4927 1094 -4853 1103
rect -4444 1094 -4370 1103
rect -4927 1038 -4918 1094
rect -4444 1038 -4435 1094
rect -4927 1029 -4853 1038
rect -4444 1029 -4370 1038
<< locali >>
rect -4648 1400 -4520 1415
rect -4648 1302 -4633 1400
rect -4535 1302 -4520 1400
rect -4304 1400 -4240 1415
rect -4648 1287 -4520 1302
rect -4439 1331 -4375 1346
rect -4439 1297 -4424 1331
rect -4390 1297 -4375 1331
rect -4439 1282 -4375 1297
rect -4304 1302 -4289 1400
rect -4255 1302 -4240 1400
rect -4304 1287 -4240 1302
rect -3568 1284 -3510 1296
rect -3568 1250 -3556 1284
rect -3522 1250 -3510 1284
rect -3568 1238 -3510 1250
rect -3724 1142 -3596 1157
rect -3724 1044 -3709 1142
rect -3611 1044 -3596 1142
rect -3456 1142 -3392 1157
rect -3724 1029 -3596 1044
rect -3555 1078 -3491 1093
rect -3555 1044 -3540 1078
rect -3506 1044 -3491 1078
rect -3555 1029 -3491 1044
rect -3456 1044 -3441 1142
rect -3407 1044 -3392 1142
rect -3456 1029 -3392 1044
rect -3610 774 -3482 789
rect -3610 740 -3595 774
rect -3497 740 -3482 774
rect -3610 725 -3482 740
rect -7515 -3410 -7451 -3395
rect -7515 -3508 -7500 -3410
rect -7466 -3508 -7451 -3410
rect -7515 -3523 -7451 -3508
rect -5403 -3410 -5339 -3395
rect -5403 -3508 -5388 -3410
rect -5354 -3508 -5339 -3410
rect -5403 -3523 -5339 -3508
rect -3291 -3410 -3227 -3395
rect -3291 -3508 -3276 -3410
rect -3242 -3508 -3227 -3410
rect -3291 -3523 -3227 -3508
rect -1179 -3410 -1115 -3395
rect -1179 -3508 -1164 -3410
rect -1130 -3508 -1115 -3410
rect -1179 -3523 -1115 -3508
rect 933 -3410 997 -3395
rect 933 -3508 948 -3410
rect 982 -3508 997 -3410
rect 933 -3523 997 -3508
rect 3045 -3410 3109 -3395
rect 3045 -3508 3060 -3410
rect 3094 -3508 3109 -3410
rect 3045 -3523 3109 -3508
rect 5157 -3410 5221 -3395
rect 5157 -3508 5172 -3410
rect 5206 -3508 5221 -3410
rect 5157 -3523 5221 -3508
rect 7269 -3410 7333 -3395
rect 7269 -3508 7284 -3410
rect 7318 -3508 7333 -3410
rect 7269 -3523 7333 -3508
rect 9381 -3410 9445 -3395
rect 9381 -3508 9396 -3410
rect 9430 -3508 9445 -3410
rect 9381 -3523 9445 -3508
rect -9047 -4142 -8983 -4127
rect -9047 -4240 -9032 -4142
rect -8998 -4240 -8983 -4142
rect -9047 -4255 -8983 -4240
rect -6935 -4142 -6871 -4127
rect -6935 -4240 -6920 -4142
rect -6886 -4240 -6871 -4142
rect -6935 -4255 -6871 -4240
rect -4823 -4142 -4759 -4127
rect -4823 -4240 -4808 -4142
rect -4774 -4240 -4759 -4142
rect -4823 -4255 -4759 -4240
rect -2711 -4142 -2647 -4127
rect -2711 -4240 -2696 -4142
rect -2662 -4240 -2647 -4142
rect -2711 -4255 -2647 -4240
rect -599 -4142 -535 -4127
rect -599 -4240 -584 -4142
rect -550 -4240 -535 -4142
rect -599 -4255 -535 -4240
rect 1513 -4142 1577 -4127
rect 1513 -4240 1528 -4142
rect 1562 -4240 1577 -4142
rect 1513 -4255 1577 -4240
rect 3625 -4142 3689 -4127
rect 3625 -4240 3640 -4142
rect 3674 -4240 3689 -4142
rect 3625 -4255 3689 -4240
rect 5737 -4142 5801 -4127
rect 5737 -4240 5752 -4142
rect 5786 -4240 5801 -4142
rect 5737 -4255 5801 -4240
rect 7849 -4142 7913 -4127
rect 7849 -4240 7864 -4142
rect 7898 -4240 7913 -4142
rect 7849 -4255 7913 -4240
rect -7515 -5144 -7451 -5129
rect -7515 -5242 -7500 -5144
rect -7466 -5242 -7451 -5144
rect -7515 -5257 -7451 -5242
rect -5403 -5144 -5339 -5129
rect -5403 -5242 -5388 -5144
rect -5354 -5242 -5339 -5144
rect -5403 -5257 -5339 -5242
rect -3291 -5144 -3227 -5129
rect -3291 -5242 -3276 -5144
rect -3242 -5242 -3227 -5144
rect -3291 -5257 -3227 -5242
rect -1179 -5144 -1115 -5129
rect -1179 -5242 -1164 -5144
rect -1130 -5242 -1115 -5144
rect -1179 -5257 -1115 -5242
rect 933 -5144 997 -5129
rect 933 -5242 948 -5144
rect 982 -5242 997 -5144
rect 933 -5257 997 -5242
rect 3045 -5144 3109 -5129
rect 3045 -5242 3060 -5144
rect 3094 -5242 3109 -5144
rect 3045 -5257 3109 -5242
rect 5157 -5144 5221 -5129
rect 5157 -5242 5172 -5144
rect 5206 -5242 5221 -5144
rect 5157 -5257 5221 -5242
rect 7269 -5144 7333 -5129
rect 7269 -5242 7284 -5144
rect 7318 -5242 7333 -5144
rect 7269 -5257 7333 -5242
rect 9381 -5144 9445 -5129
rect 9381 -5242 9396 -5144
rect 9430 -5242 9445 -5144
rect 9381 -5257 9445 -5242
rect -9047 -5876 -8983 -5861
rect -9047 -5974 -9032 -5876
rect -8998 -5974 -8983 -5876
rect -9047 -5989 -8983 -5974
rect -6935 -5876 -6871 -5861
rect -6935 -5974 -6920 -5876
rect -6886 -5974 -6871 -5876
rect -6935 -5989 -6871 -5974
rect -4823 -5876 -4759 -5861
rect -4823 -5974 -4808 -5876
rect -4774 -5974 -4759 -5876
rect -4823 -5989 -4759 -5974
rect -2711 -5876 -2647 -5861
rect -2711 -5974 -2696 -5876
rect -2662 -5974 -2647 -5876
rect -2711 -5989 -2647 -5974
rect -599 -5876 -535 -5861
rect -599 -5974 -584 -5876
rect -550 -5974 -535 -5876
rect -599 -5989 -535 -5974
rect 1513 -5876 1577 -5861
rect 1513 -5974 1528 -5876
rect 1562 -5974 1577 -5876
rect 1513 -5989 1577 -5974
rect 3625 -5876 3689 -5861
rect 3625 -5974 3640 -5876
rect 3674 -5974 3689 -5876
rect 3625 -5989 3689 -5974
rect 5737 -5876 5801 -5861
rect 5737 -5974 5752 -5876
rect 5786 -5974 5801 -5876
rect 5737 -5989 5801 -5974
rect 7849 -5876 7913 -5861
rect 7849 -5974 7864 -5876
rect 7898 -5974 7913 -5876
rect 7849 -5989 7913 -5974
<< viali >>
rect -4633 1302 -4535 1400
rect -4424 1297 -4390 1331
rect -4289 1302 -4255 1400
rect -3556 1250 -3522 1284
rect -3709 1044 -3611 1142
rect -3540 1044 -3506 1078
rect -3441 1044 -3407 1142
rect -3595 740 -3497 774
rect -7500 -3508 -7466 -3410
rect -5388 -3508 -5354 -3410
rect -3276 -3508 -3242 -3410
rect -1164 -3508 -1130 -3410
rect 948 -3508 982 -3410
rect 3060 -3508 3094 -3410
rect 5172 -3508 5206 -3410
rect 7284 -3508 7318 -3410
rect 9396 -3508 9430 -3410
rect -9032 -4240 -8998 -4142
rect -6920 -4240 -6886 -4142
rect -4808 -4240 -4774 -4142
rect -2696 -4240 -2662 -4142
rect -584 -4240 -550 -4142
rect 1528 -4240 1562 -4142
rect 3640 -4240 3674 -4142
rect 5752 -4240 5786 -4142
rect 7864 -4240 7898 -4142
rect -7500 -5242 -7466 -5144
rect -5388 -5242 -5354 -5144
rect -3276 -5242 -3242 -5144
rect -1164 -5242 -1130 -5144
rect 948 -5242 982 -5144
rect 3060 -5242 3094 -5144
rect 5172 -5242 5206 -5144
rect 7284 -5242 7318 -5144
rect 9396 -5242 9430 -5144
rect -9032 -5974 -8998 -5876
rect -6920 -5974 -6886 -5876
rect -4808 -5974 -4774 -5876
rect -2696 -5974 -2662 -5876
rect -584 -5974 -550 -5876
rect 1528 -5974 1562 -5876
rect 3640 -5974 3674 -5876
rect 5752 -5974 5786 -5876
rect 7864 -5974 7898 -5876
<< metal1 >>
rect -4658 1414 -4510 1425
rect -4658 1288 -4647 1414
rect -4521 1288 -4510 1414
rect -4309 1414 -4235 1425
rect -4658 1277 -4510 1288
rect -4444 1340 -4370 1351
rect -4444 1288 -4433 1340
rect -4381 1288 -4370 1340
rect -4444 1277 -4370 1288
rect -4309 1288 -4298 1414
rect -4246 1288 -4235 1414
rect -4309 1277 -4235 1288
rect -3568 1284 -3510 1296
rect -3568 1250 -3556 1284
rect -3522 1250 -3510 1284
rect -3568 1238 -3510 1250
rect -4658 1166 -4510 1177
rect -4658 1040 -4647 1166
rect -4521 1040 -4510 1166
rect -4309 1166 -4235 1177
rect -4658 1029 -4510 1040
rect -4444 1092 -4370 1103
rect -4444 1040 -4433 1092
rect -4381 1040 -4370 1092
rect -4444 1029 -4370 1040
rect -4309 1040 -4298 1166
rect -4246 1040 -4235 1166
rect -4309 1029 -4235 1040
rect -4152 1151 -4024 1157
rect -4152 1035 -4146 1151
rect -4030 1035 -4024 1151
rect -3884 1151 -3820 1157
rect -4152 1029 -4024 1035
rect -3983 1087 -3919 1093
rect -3983 1035 -3977 1087
rect -3925 1035 -3919 1087
rect -3983 1029 -3919 1035
rect -3884 1035 -3878 1151
rect -3826 1035 -3820 1151
rect -3884 1029 -3820 1035
rect -3724 1151 -3596 1157
rect -3724 1035 -3718 1151
rect -3602 1035 -3596 1151
rect -3456 1151 -3392 1157
rect -3724 1029 -3596 1035
rect -3555 1087 -3491 1093
rect -3555 1035 -3549 1087
rect -3497 1035 -3491 1087
rect -3555 1029 -3491 1035
rect -3456 1035 -3450 1151
rect -3398 1035 -3392 1151
rect -3456 1029 -3392 1035
rect -3864 857 -3736 863
rect -3864 805 -3858 857
rect -3742 805 -3736 857
rect -3864 799 -3736 805
rect -3610 783 -3482 789
rect -4300 768 -4152 779
rect -4300 716 -4289 768
rect -4163 716 -4152 768
rect -3610 731 -3604 783
rect -3488 731 -3482 783
rect -3610 725 -3482 731
rect -4300 705 -4152 716
rect -9852 -2918 9468 -2912
rect -9852 -3054 -9846 -2918
rect -9730 -3054 9468 -2918
rect -9852 -3060 9468 -3054
rect -7515 -3401 -7451 -3395
rect -7515 -3517 -7509 -3401
rect -7457 -3517 -7451 -3401
rect -7515 -3523 -7451 -3517
rect -5403 -3401 -5339 -3395
rect -5403 -3517 -5397 -3401
rect -5345 -3517 -5339 -3401
rect -5403 -3523 -5339 -3517
rect -3291 -3401 -3227 -3395
rect -3291 -3517 -3285 -3401
rect -3233 -3517 -3227 -3401
rect -3291 -3523 -3227 -3517
rect -1179 -3401 -1115 -3395
rect -1179 -3517 -1173 -3401
rect -1121 -3517 -1115 -3401
rect -1179 -3523 -1115 -3517
rect 933 -3401 997 -3395
rect 933 -3517 939 -3401
rect 991 -3517 997 -3401
rect 933 -3523 997 -3517
rect 3045 -3401 3109 -3395
rect 3045 -3517 3051 -3401
rect 3103 -3517 3109 -3401
rect 3045 -3523 3109 -3517
rect 5157 -3401 5221 -3395
rect 5157 -3517 5163 -3401
rect 5215 -3517 5221 -3401
rect 5157 -3523 5221 -3517
rect 7269 -3401 7333 -3395
rect 7269 -3517 7275 -3401
rect 7327 -3517 7333 -3401
rect 7269 -3523 7333 -3517
rect 9381 -3401 9445 -3395
rect 9381 -3517 9387 -3401
rect 9439 -3517 9445 -3401
rect 9381 -3523 9445 -3517
rect -10052 -3630 9468 -3624
rect -10052 -3868 -10046 -3630
rect -9930 -3868 9468 -3630
rect -10052 -3874 9468 -3868
rect -10252 -3904 -9526 -3902
rect -10252 -3956 -10246 -3904
rect -10130 -3956 -9526 -3904
rect -10252 -3959 -9526 -3956
rect -7442 -3959 -7414 -3902
rect -5330 -3959 -5302 -3902
rect -3218 -3959 -3190 -3902
rect -1106 -3959 -1078 -3902
rect 1006 -3959 1034 -3902
rect 3118 -3959 3146 -3902
rect 5230 -3959 5258 -3902
rect 7342 -3959 7370 -3902
rect 9454 -3959 9468 -3902
rect -9047 -4133 -8983 -4127
rect -9047 -4249 -9041 -4133
rect -8989 -4249 -8983 -4133
rect -9047 -4255 -8983 -4249
rect -6935 -4133 -6871 -4127
rect -6935 -4249 -6929 -4133
rect -6877 -4249 -6871 -4133
rect -6935 -4255 -6871 -4249
rect -4823 -4133 -4759 -4127
rect -4823 -4249 -4817 -4133
rect -4765 -4249 -4759 -4133
rect -4823 -4255 -4759 -4249
rect -2711 -4133 -2647 -4127
rect -2711 -4249 -2705 -4133
rect -2653 -4249 -2647 -4133
rect -2711 -4255 -2647 -4249
rect -599 -4133 -535 -4127
rect -599 -4249 -593 -4133
rect -541 -4249 -535 -4133
rect -599 -4255 -535 -4249
rect 1513 -4133 1577 -4127
rect 1513 -4249 1519 -4133
rect 1571 -4249 1577 -4133
rect 1513 -4255 1577 -4249
rect 3625 -4133 3689 -4127
rect 3625 -4249 3631 -4133
rect 3683 -4249 3689 -4133
rect 3625 -4255 3689 -4249
rect 5737 -4133 5801 -4127
rect 5737 -4249 5743 -4133
rect 5795 -4249 5801 -4133
rect 5737 -4255 5801 -4249
rect 7849 -4133 7913 -4127
rect 7849 -4249 7855 -4133
rect 7907 -4249 7913 -4133
rect 7849 -4255 7913 -4249
rect -9852 -4444 9468 -4438
rect -9852 -4788 -9846 -4444
rect -9730 -4788 9468 -4444
rect -9852 -4794 9468 -4788
rect -7515 -5135 -7451 -5129
rect -7515 -5251 -7509 -5135
rect -7457 -5251 -7451 -5135
rect -7515 -5257 -7451 -5251
rect -5403 -5135 -5339 -5129
rect -5403 -5251 -5397 -5135
rect -5345 -5251 -5339 -5135
rect -5403 -5257 -5339 -5251
rect -3291 -5135 -3227 -5129
rect -3291 -5251 -3285 -5135
rect -3233 -5251 -3227 -5135
rect -3291 -5257 -3227 -5251
rect -1179 -5135 -1115 -5129
rect -1179 -5251 -1173 -5135
rect -1121 -5251 -1115 -5135
rect -1179 -5257 -1115 -5251
rect 933 -5135 997 -5129
rect 933 -5251 939 -5135
rect 991 -5251 997 -5135
rect 933 -5257 997 -5251
rect 3045 -5135 3109 -5129
rect 3045 -5251 3051 -5135
rect 3103 -5251 3109 -5135
rect 3045 -5257 3109 -5251
rect 5157 -5135 5221 -5129
rect 5157 -5251 5163 -5135
rect 5215 -5251 5221 -5135
rect 5157 -5257 5221 -5251
rect 7269 -5135 7333 -5129
rect 7269 -5251 7275 -5135
rect 7327 -5251 7333 -5135
rect 7269 -5257 7333 -5251
rect 9381 -5135 9445 -5129
rect 9381 -5251 9387 -5135
rect 9439 -5251 9445 -5135
rect 9381 -5257 9445 -5251
rect -10052 -5364 9468 -5358
rect -10052 -5602 -10046 -5364
rect -9930 -5602 9468 -5364
rect -10052 -5608 9468 -5602
rect -10252 -5638 -9526 -5636
rect -10252 -5690 -10246 -5638
rect -10130 -5690 -9526 -5638
rect -10252 -5693 -9526 -5690
rect -7442 -5693 -7414 -5636
rect -5330 -5693 -5302 -5636
rect -3218 -5693 -3190 -5636
rect -1106 -5693 -1078 -5636
rect 1006 -5693 1034 -5636
rect 3118 -5693 3146 -5636
rect 5230 -5693 5258 -5636
rect 7342 -5693 7370 -5636
rect 9454 -5693 9468 -5636
rect -9047 -5867 -8983 -5861
rect -9047 -5983 -9041 -5867
rect -8989 -5983 -8983 -5867
rect -9047 -5989 -8983 -5983
rect -6935 -5867 -6871 -5861
rect -6935 -5983 -6929 -5867
rect -6877 -5983 -6871 -5867
rect -6935 -5989 -6871 -5983
rect -4823 -5867 -4759 -5861
rect -4823 -5983 -4817 -5867
rect -4765 -5983 -4759 -5867
rect -4823 -5989 -4759 -5983
rect -2711 -5867 -2647 -5861
rect -2711 -5983 -2705 -5867
rect -2653 -5983 -2647 -5867
rect -2711 -5989 -2647 -5983
rect -599 -5867 -535 -5861
rect -599 -5983 -593 -5867
rect -541 -5983 -535 -5867
rect -599 -5989 -535 -5983
rect 1513 -5867 1577 -5861
rect 1513 -5983 1519 -5867
rect 1571 -5983 1577 -5867
rect 1513 -5989 1577 -5983
rect 3625 -5867 3689 -5861
rect 3625 -5983 3631 -5867
rect 3683 -5983 3689 -5867
rect 3625 -5989 3689 -5983
rect 5737 -5867 5801 -5861
rect 5737 -5983 5743 -5867
rect 5795 -5983 5801 -5867
rect 5737 -5989 5801 -5983
rect 7849 -5867 7913 -5861
rect 7849 -5983 7855 -5867
rect 7907 -5983 7913 -5867
rect 7849 -5989 7913 -5983
rect -9852 -6178 9468 -6172
rect -9852 -6282 -9846 -6178
rect -10252 -6314 -9846 -6282
rect -9730 -6288 9468 -6178
rect -9730 -6314 -4574 -6288
rect -10252 -6476 -4574 -6314
rect -4386 -6476 9468 -6288
rect -10252 -6482 9468 -6476
rect -10252 -6544 9468 -6538
rect -10252 -6732 -10246 -6544
rect -10130 -6732 9468 -6544
rect -10252 -6738 9468 -6732
rect -10252 -6800 9468 -6794
rect -10252 -6988 -10046 -6800
rect -9930 -6988 9468 -6800
rect -10252 -6994 9468 -6988
rect -27806 -10519 -27406 -10513
rect -27806 -10796 -27800 -10519
rect -27412 -10796 -27406 -10519
rect -27806 -10802 -27406 -10796
rect -19274 -10802 -10164 -10552
rect -10355 -10824 -10164 -10802
rect -10355 -10830 -4887 -10824
rect -28262 -10858 -27459 -10852
rect -28262 -11096 -28256 -10858
rect -27868 -11096 -27459 -10858
rect -28262 -11102 -27459 -11096
rect -19020 -11080 -10420 -10854
rect -10355 -11018 -5076 -10830
rect -4893 -11018 -4887 -10830
rect -10355 -11024 -4887 -11018
rect -19020 -11104 -4637 -11080
rect -10614 -11280 -4637 -11104
<< via1 >>
rect -4647 1400 -4521 1414
rect -4647 1302 -4633 1400
rect -4633 1302 -4535 1400
rect -4535 1302 -4521 1400
rect -4647 1288 -4521 1302
rect -4433 1331 -4381 1340
rect -4433 1297 -4424 1331
rect -4424 1297 -4390 1331
rect -4390 1297 -4381 1331
rect -4433 1288 -4381 1297
rect -4298 1400 -4246 1414
rect -4298 1302 -4289 1400
rect -4289 1302 -4255 1400
rect -4255 1302 -4246 1400
rect -4298 1288 -4246 1302
rect -4647 1040 -4521 1166
rect -4433 1040 -4381 1092
rect -4298 1040 -4246 1166
rect -4146 1035 -4030 1151
rect -3977 1035 -3925 1087
rect -3878 1035 -3826 1151
rect -3718 1142 -3602 1151
rect -3718 1044 -3709 1142
rect -3709 1044 -3611 1142
rect -3611 1044 -3602 1142
rect -3718 1035 -3602 1044
rect -3549 1078 -3497 1087
rect -3549 1044 -3540 1078
rect -3540 1044 -3506 1078
rect -3506 1044 -3497 1078
rect -3549 1035 -3497 1044
rect -3450 1142 -3398 1151
rect -3450 1044 -3441 1142
rect -3441 1044 -3407 1142
rect -3407 1044 -3398 1142
rect -3450 1035 -3398 1044
rect -3858 805 -3742 857
rect -4289 716 -4163 768
rect -3604 774 -3488 783
rect -3604 740 -3595 774
rect -3595 740 -3497 774
rect -3497 740 -3488 774
rect -3604 731 -3488 740
rect -9846 -3054 -9730 -2918
rect -7509 -3410 -7457 -3401
rect -7509 -3508 -7500 -3410
rect -7500 -3508 -7466 -3410
rect -7466 -3508 -7457 -3410
rect -7509 -3517 -7457 -3508
rect -5397 -3410 -5345 -3401
rect -5397 -3508 -5388 -3410
rect -5388 -3508 -5354 -3410
rect -5354 -3508 -5345 -3410
rect -5397 -3517 -5345 -3508
rect -3285 -3410 -3233 -3401
rect -3285 -3508 -3276 -3410
rect -3276 -3508 -3242 -3410
rect -3242 -3508 -3233 -3410
rect -3285 -3517 -3233 -3508
rect -1173 -3410 -1121 -3401
rect -1173 -3508 -1164 -3410
rect -1164 -3508 -1130 -3410
rect -1130 -3508 -1121 -3410
rect -1173 -3517 -1121 -3508
rect 939 -3410 991 -3401
rect 939 -3508 948 -3410
rect 948 -3508 982 -3410
rect 982 -3508 991 -3410
rect 939 -3517 991 -3508
rect 3051 -3410 3103 -3401
rect 3051 -3508 3060 -3410
rect 3060 -3508 3094 -3410
rect 3094 -3508 3103 -3410
rect 3051 -3517 3103 -3508
rect 5163 -3410 5215 -3401
rect 5163 -3508 5172 -3410
rect 5172 -3508 5206 -3410
rect 5206 -3508 5215 -3410
rect 5163 -3517 5215 -3508
rect 7275 -3410 7327 -3401
rect 7275 -3508 7284 -3410
rect 7284 -3508 7318 -3410
rect 7318 -3508 7327 -3410
rect 7275 -3517 7327 -3508
rect 9387 -3410 9439 -3401
rect 9387 -3508 9396 -3410
rect 9396 -3508 9430 -3410
rect 9430 -3508 9439 -3410
rect 9387 -3517 9439 -3508
rect -10046 -3868 -9930 -3630
rect -10246 -3956 -10130 -3904
rect -9041 -4142 -8989 -4133
rect -9041 -4240 -9032 -4142
rect -9032 -4240 -8998 -4142
rect -8998 -4240 -8989 -4142
rect -9041 -4249 -8989 -4240
rect -6929 -4142 -6877 -4133
rect -6929 -4240 -6920 -4142
rect -6920 -4240 -6886 -4142
rect -6886 -4240 -6877 -4142
rect -6929 -4249 -6877 -4240
rect -4817 -4142 -4765 -4133
rect -4817 -4240 -4808 -4142
rect -4808 -4240 -4774 -4142
rect -4774 -4240 -4765 -4142
rect -4817 -4249 -4765 -4240
rect -2705 -4142 -2653 -4133
rect -2705 -4240 -2696 -4142
rect -2696 -4240 -2662 -4142
rect -2662 -4240 -2653 -4142
rect -2705 -4249 -2653 -4240
rect -593 -4142 -541 -4133
rect -593 -4240 -584 -4142
rect -584 -4240 -550 -4142
rect -550 -4240 -541 -4142
rect -593 -4249 -541 -4240
rect 1519 -4142 1571 -4133
rect 1519 -4240 1528 -4142
rect 1528 -4240 1562 -4142
rect 1562 -4240 1571 -4142
rect 1519 -4249 1571 -4240
rect 3631 -4142 3683 -4133
rect 3631 -4240 3640 -4142
rect 3640 -4240 3674 -4142
rect 3674 -4240 3683 -4142
rect 3631 -4249 3683 -4240
rect 5743 -4142 5795 -4133
rect 5743 -4240 5752 -4142
rect 5752 -4240 5786 -4142
rect 5786 -4240 5795 -4142
rect 5743 -4249 5795 -4240
rect 7855 -4142 7907 -4133
rect 7855 -4240 7864 -4142
rect 7864 -4240 7898 -4142
rect 7898 -4240 7907 -4142
rect 7855 -4249 7907 -4240
rect -9846 -4788 -9730 -4444
rect -7509 -5144 -7457 -5135
rect -7509 -5242 -7500 -5144
rect -7500 -5242 -7466 -5144
rect -7466 -5242 -7457 -5144
rect -7509 -5251 -7457 -5242
rect -5397 -5144 -5345 -5135
rect -5397 -5242 -5388 -5144
rect -5388 -5242 -5354 -5144
rect -5354 -5242 -5345 -5144
rect -5397 -5251 -5345 -5242
rect -3285 -5144 -3233 -5135
rect -3285 -5242 -3276 -5144
rect -3276 -5242 -3242 -5144
rect -3242 -5242 -3233 -5144
rect -3285 -5251 -3233 -5242
rect -1173 -5144 -1121 -5135
rect -1173 -5242 -1164 -5144
rect -1164 -5242 -1130 -5144
rect -1130 -5242 -1121 -5144
rect -1173 -5251 -1121 -5242
rect 939 -5144 991 -5135
rect 939 -5242 948 -5144
rect 948 -5242 982 -5144
rect 982 -5242 991 -5144
rect 939 -5251 991 -5242
rect 3051 -5144 3103 -5135
rect 3051 -5242 3060 -5144
rect 3060 -5242 3094 -5144
rect 3094 -5242 3103 -5144
rect 3051 -5251 3103 -5242
rect 5163 -5144 5215 -5135
rect 5163 -5242 5172 -5144
rect 5172 -5242 5206 -5144
rect 5206 -5242 5215 -5144
rect 5163 -5251 5215 -5242
rect 7275 -5144 7327 -5135
rect 7275 -5242 7284 -5144
rect 7284 -5242 7318 -5144
rect 7318 -5242 7327 -5144
rect 7275 -5251 7327 -5242
rect 9387 -5144 9439 -5135
rect 9387 -5242 9396 -5144
rect 9396 -5242 9430 -5144
rect 9430 -5242 9439 -5144
rect 9387 -5251 9439 -5242
rect -10046 -5602 -9930 -5364
rect -10246 -5690 -10130 -5638
rect -9041 -5876 -8989 -5867
rect -9041 -5974 -9032 -5876
rect -9032 -5974 -8998 -5876
rect -8998 -5974 -8989 -5876
rect -9041 -5983 -8989 -5974
rect -6929 -5876 -6877 -5867
rect -6929 -5974 -6920 -5876
rect -6920 -5974 -6886 -5876
rect -6886 -5974 -6877 -5876
rect -6929 -5983 -6877 -5974
rect -4817 -5876 -4765 -5867
rect -4817 -5974 -4808 -5876
rect -4808 -5974 -4774 -5876
rect -4774 -5974 -4765 -5876
rect -4817 -5983 -4765 -5974
rect -2705 -5876 -2653 -5867
rect -2705 -5974 -2696 -5876
rect -2696 -5974 -2662 -5876
rect -2662 -5974 -2653 -5876
rect -2705 -5983 -2653 -5974
rect -593 -5876 -541 -5867
rect -593 -5974 -584 -5876
rect -584 -5974 -550 -5876
rect -550 -5974 -541 -5876
rect -593 -5983 -541 -5974
rect 1519 -5876 1571 -5867
rect 1519 -5974 1528 -5876
rect 1528 -5974 1562 -5876
rect 1562 -5974 1571 -5876
rect 1519 -5983 1571 -5974
rect 3631 -5876 3683 -5867
rect 3631 -5974 3640 -5876
rect 3640 -5974 3674 -5876
rect 3674 -5974 3683 -5876
rect 3631 -5983 3683 -5974
rect 5743 -5876 5795 -5867
rect 5743 -5974 5752 -5876
rect 5752 -5974 5786 -5876
rect 5786 -5974 5795 -5876
rect 5743 -5983 5795 -5974
rect 7855 -5876 7907 -5867
rect 7855 -5974 7864 -5876
rect 7864 -5974 7898 -5876
rect 7898 -5974 7907 -5876
rect 7855 -5983 7907 -5974
rect -9846 -6314 -9730 -6178
rect -4574 -6476 -4386 -6288
rect -10246 -6732 -10130 -6544
rect -10046 -6988 -9930 -6800
rect -4574 -7700 -4386 -7564
rect -27800 -10796 -27412 -10519
rect -28256 -11096 -27868 -10858
rect -5076 -11018 -4893 -10830
rect -4575 -11018 -4387 -10830
<< metal2 >>
rect -28262 10255 -27862 10398
rect -28262 10119 -27929 10255
rect -27868 10119 -27862 10255
rect -28262 -10858 -27862 10119
rect -27806 6812 -27406 10398
rect -19249 7756 -19185 7760
rect -19254 7751 -19180 7756
rect -19254 7687 -19249 7751
rect -19185 7687 -19180 7751
rect -27035 7147 -26979 7156
rect -27035 7082 -26979 7091
rect -27806 6676 -27478 6812
rect -27412 6676 -27406 6812
rect -27806 2314 -27406 6676
rect -27806 2178 -27478 2314
rect -27412 2178 -27406 2314
rect -27806 -10519 -27406 2178
rect -19254 607 -19180 7687
rect -17661 7151 -17597 7160
rect -18588 5514 -18528 5523
rect -18588 -8044 -18528 5454
rect -18293 5314 -18229 5323
rect -18293 2438 -18229 5250
rect -18293 2374 -18177 2438
rect -18241 -2878 -18177 2374
rect -17661 -2678 -17597 7087
rect -4658 1416 -4510 1425
rect -4658 1286 -4649 1416
rect -4519 1286 -4510 1416
rect -4309 1416 -4235 1425
rect -4658 1277 -4510 1286
rect -4444 1342 -4370 1351
rect -4444 1286 -4435 1342
rect -4379 1286 -4370 1342
rect -4444 1277 -4370 1286
rect -4309 1286 -4300 1416
rect -4244 1286 -4235 1416
rect -4309 1277 -4235 1286
rect -5142 1168 -4994 1177
rect -5142 1038 -5133 1168
rect -5003 1038 -4994 1168
rect -4793 1168 -4719 1177
rect -5142 1029 -4994 1038
rect -4927 1094 -4853 1103
rect -4927 1038 -4918 1094
rect -4862 1038 -4853 1094
rect -4927 1029 -4853 1038
rect -4793 1038 -4784 1168
rect -4728 1038 -4719 1168
rect -4793 1029 -4719 1038
rect -4658 1168 -4510 1177
rect -4658 1038 -4649 1168
rect -4519 1038 -4510 1168
rect -4309 1168 -4235 1177
rect -4658 1029 -4510 1038
rect -4444 1094 -4370 1103
rect -4444 1038 -4435 1094
rect -4379 1038 -4370 1094
rect -4444 1029 -4370 1038
rect -4309 1038 -4300 1168
rect -4244 1038 -4235 1168
rect -4309 1029 -4235 1038
rect -4152 1151 -4024 1157
rect -4152 1035 -4146 1151
rect -4030 1035 -4024 1151
rect -3884 1151 -3820 1157
rect -4152 1029 -4024 1035
rect -3983 1087 -3919 1093
rect -3983 1035 -3977 1087
rect -3925 1035 -3919 1087
rect -3983 1029 -3919 1035
rect -3884 1035 -3878 1151
rect -3826 1035 -3820 1151
rect -3884 1029 -3820 1035
rect -3724 1151 -3596 1157
rect -3724 1035 -3718 1151
rect -3602 1035 -3596 1151
rect -3456 1151 -3392 1157
rect -3724 1029 -3596 1035
rect -3555 1087 -3491 1093
rect -3555 1035 -3549 1087
rect -3497 1035 -3491 1087
rect -3555 1029 -3491 1035
rect -3456 1035 -3450 1151
rect -3398 1035 -3392 1151
rect -3456 1029 -3392 1035
rect -3864 857 -3736 863
rect -4784 814 -4636 823
rect -4784 758 -4775 814
rect -4645 758 -4636 814
rect -3864 805 -3858 857
rect -3742 805 -3736 857
rect -3864 799 -3736 805
rect -3610 783 -3482 789
rect -17531 605 -17457 753
rect -4784 749 -4636 758
rect -4300 770 -4152 779
rect -4300 714 -4291 770
rect -4161 714 -4152 770
rect -3610 731 -3604 783
rect -3488 731 -3482 783
rect -3610 725 -3482 731
rect -4300 705 -4152 714
rect -12959 -903 -12895 -894
rect -15351 -2196 -15287 -2068
rect -17666 -2734 -17657 -2678
rect -17601 -2734 -17592 -2678
rect -17661 -2738 -17597 -2734
rect -13162 -2745 -13084 -2709
rect -13162 -7524 -13098 -2745
rect -12959 -3378 -12895 -967
rect -12959 -3434 -12955 -3378
rect -12899 -3434 -12895 -3378
rect -12959 -3438 -12895 -3434
rect -12955 -3443 -12899 -3438
rect -10252 -3904 -10124 -2912
rect -10252 -3956 -10246 -3904
rect -10130 -3956 -10124 -3904
rect -10252 -5638 -10124 -3956
rect -10252 -5690 -10246 -5638
rect -10130 -5690 -10124 -5638
rect -10252 -6544 -10124 -5690
rect -10252 -6732 -10246 -6544
rect -10130 -6732 -10124 -6544
rect -10252 -6738 -10124 -6732
rect -10052 -3630 -9924 -2912
rect -10052 -3868 -10046 -3630
rect -9930 -3868 -9924 -3630
rect -10052 -5364 -9924 -3868
rect -10052 -5602 -10046 -5364
rect -9930 -5602 -9924 -5364
rect -10052 -6800 -9924 -5602
rect -9852 -2918 -9724 -2912
rect -9852 -3054 -9846 -2918
rect -9730 -3054 -9724 -2918
rect -9852 -4444 -9724 -3054
rect -9597 -3374 -9533 -3365
rect -9597 -3690 -9533 -3438
rect -7515 -3401 -7451 -3395
rect -7515 -3517 -7509 -3401
rect -7457 -3517 -7451 -3401
rect -9602 -3746 -9593 -3690
rect -9537 -3746 -9528 -3690
rect -9597 -3750 -9533 -3746
rect -9047 -4133 -8983 -4127
rect -9047 -4249 -9041 -4133
rect -8989 -4249 -8983 -4133
rect -9047 -4319 -8983 -4249
rect -9852 -4788 -9846 -4444
rect -9730 -4788 -9724 -4444
rect -9852 -6178 -9724 -4788
rect -7515 -4996 -7451 -3517
rect -5403 -3401 -5339 -3395
rect -5403 -3517 -5397 -3401
rect -5345 -3517 -5339 -3401
rect -6935 -4133 -6871 -4127
rect -6935 -4249 -6929 -4133
rect -6877 -4249 -6871 -4133
rect -6935 -4319 -6871 -4249
rect -5403 -4967 -5339 -3517
rect -3291 -3401 -3227 -3395
rect -3291 -3517 -3285 -3401
rect -3233 -3517 -3227 -3401
rect -4823 -4133 -4759 -4127
rect -4823 -4249 -4817 -4133
rect -4765 -4249 -4759 -4133
rect -4823 -4319 -4759 -4249
rect -3291 -4945 -3227 -3517
rect -1179 -3401 -1115 -3395
rect -1179 -3517 -1173 -3401
rect -1121 -3517 -1115 -3401
rect -2711 -4133 -2647 -4127
rect -2711 -4249 -2705 -4133
rect -2653 -4249 -2647 -4133
rect -2711 -4319 -2647 -4249
rect -1179 -4924 -1115 -3517
rect 933 -3401 997 -3395
rect 933 -3517 939 -3401
rect 991 -3517 997 -3401
rect -599 -4133 -535 -4127
rect -599 -4249 -593 -4133
rect -541 -4249 -535 -4133
rect -599 -4319 -535 -4249
rect -7515 -5060 -7341 -4996
rect -5403 -5031 -5223 -4967
rect -3291 -5009 -3111 -4945
rect -1179 -4988 -956 -4924
rect -7515 -5135 -7451 -5129
rect -7515 -5251 -7509 -5135
rect -7457 -5251 -7451 -5135
rect -9047 -5867 -8983 -5861
rect -9047 -5983 -9041 -5867
rect -8989 -5983 -8983 -5867
rect -9047 -6053 -8983 -5983
rect -9852 -6314 -9846 -6178
rect -9730 -6314 -9724 -6178
rect -9852 -6320 -9724 -6314
rect -10052 -6988 -10046 -6800
rect -9930 -6988 -9924 -6800
rect -10052 -6994 -9924 -6988
rect -7515 -7298 -7451 -5251
rect -7405 -7152 -7341 -5060
rect -5403 -5135 -5339 -5129
rect -5403 -5251 -5397 -5135
rect -5345 -5251 -5339 -5135
rect -6935 -5867 -6871 -5861
rect -6935 -5983 -6929 -5867
rect -6877 -5983 -6871 -5867
rect -6935 -6053 -6871 -5983
rect -5403 -7014 -5339 -5251
rect -5287 -6876 -5223 -5031
rect -3291 -5135 -3227 -5129
rect -3291 -5251 -3285 -5135
rect -3233 -5251 -3227 -5135
rect -4823 -5867 -4759 -5861
rect -4823 -5983 -4817 -5867
rect -4765 -5983 -4759 -5867
rect -4823 -6053 -4759 -5983
rect -5287 -6949 -5223 -6940
rect -4580 -6288 -4380 -6282
rect -4580 -6476 -4574 -6288
rect -4386 -6476 -4380 -6288
rect -5403 -7087 -5339 -7078
rect -7405 -7225 -7341 -7216
rect -7515 -7371 -7451 -7362
rect -5084 -7520 -5028 -7515
rect -13162 -7580 -13158 -7524
rect -13102 -7580 -13098 -7524
rect -13162 -7584 -13098 -7580
rect -5088 -7524 -5024 -7520
rect -5088 -7580 -5084 -7524
rect -5028 -7580 -5024 -7524
rect -13158 -7589 -13102 -7584
rect -18588 -8100 -18586 -8044
rect -18530 -8100 -18528 -8044
rect -18588 -8102 -18528 -8100
rect -18586 -8109 -18530 -8102
rect -5088 -8780 -5024 -7580
rect -4580 -7564 -4380 -6476
rect -3291 -6710 -3227 -5251
rect -3175 -6544 -3111 -5009
rect -1179 -5135 -1115 -5129
rect -1179 -5251 -1173 -5135
rect -1121 -5251 -1115 -5135
rect -2711 -5867 -2647 -5861
rect -2711 -5983 -2705 -5867
rect -2653 -5983 -2647 -5867
rect -2711 -6053 -2647 -5983
rect -1529 -6544 -1473 -6539
rect -3175 -6617 -3111 -6608
rect -1533 -6548 -1469 -6544
rect -1533 -6604 -1529 -6548
rect -1473 -6604 -1469 -6548
rect -2079 -6710 -2023 -6705
rect -3291 -6783 -3227 -6774
rect -2083 -6714 -2019 -6710
rect -2083 -6770 -2079 -6714
rect -2023 -6770 -2019 -6714
rect -2614 -6876 -2558 -6871
rect -2618 -6880 -2554 -6876
rect -2618 -6936 -2614 -6880
rect -2558 -6936 -2554 -6880
rect -3142 -7014 -3086 -7009
rect -3146 -7018 -3082 -7014
rect -3146 -7074 -3142 -7018
rect -3086 -7074 -3082 -7018
rect -3666 -7152 -3610 -7147
rect -3670 -7156 -3606 -7152
rect -3670 -7212 -3666 -7156
rect -3610 -7212 -3606 -7156
rect -4212 -7302 -4156 -7293
rect -4212 -7367 -4156 -7358
rect -3670 -7371 -3606 -7212
rect -3146 -7382 -3082 -7074
rect -2618 -7374 -2554 -6936
rect -2083 -7374 -2019 -6770
rect -1533 -7374 -1469 -6604
rect -1179 -7303 -1115 -5251
rect -1020 -7122 -956 -4988
rect 933 -4982 997 -3517
rect 3045 -3401 3109 -3395
rect 3045 -3517 3051 -3401
rect 3103 -3517 3109 -3401
rect 1513 -4133 1577 -4127
rect 1513 -4249 1519 -4133
rect 1571 -4249 1577 -4133
rect 1513 -4319 1577 -4249
rect 3045 -4978 3109 -3517
rect 5157 -3401 5221 -3395
rect 5157 -3517 5163 -3401
rect 5215 -3517 5221 -3401
rect 3625 -4133 3689 -4127
rect 3625 -4249 3631 -4133
rect 3683 -4249 3689 -4133
rect 3625 -4319 3689 -4249
rect 5157 -4971 5221 -3517
rect 7269 -3401 7333 -3395
rect 7269 -3517 7275 -3401
rect 7327 -3517 7333 -3401
rect 5737 -4133 5801 -4127
rect 5737 -4249 5743 -4133
rect 5795 -4249 5801 -4133
rect 5737 -4319 5801 -4249
rect 7269 -4942 7333 -3517
rect 9381 -3401 9445 -3395
rect 9381 -3517 9387 -3401
rect 9439 -3517 9445 -3401
rect 9381 -3686 9445 -3517
rect 9381 -3759 9445 -3750
rect 7849 -4133 7913 -4127
rect 7849 -4249 7855 -4133
rect 7907 -4249 7913 -4133
rect 7849 -4319 7913 -4249
rect 933 -5046 1149 -4982
rect 3045 -5042 3247 -4978
rect 5157 -5035 5367 -4971
rect 7269 -5006 7480 -4942
rect 933 -5135 997 -5129
rect 933 -5251 939 -5135
rect 991 -5251 997 -5135
rect -599 -5867 -535 -5861
rect -599 -5983 -593 -5867
rect -541 -5983 -535 -5867
rect -599 -6053 -535 -5983
rect 76 -6059 132 -6054
rect 933 -6059 997 -5251
rect 72 -6063 136 -6059
rect 72 -6119 76 -6063
rect 132 -6119 136 -6063
rect -466 -7122 -410 -7117
rect -1020 -7195 -956 -7186
rect -470 -7126 -406 -7122
rect -470 -7182 -466 -7126
rect -410 -7182 -406 -7126
rect -1179 -7367 -934 -7303
rect -470 -7382 -406 -7182
rect 72 -7374 136 -6119
rect 933 -6132 997 -6123
rect 597 -6197 653 -6192
rect 1085 -6197 1149 -5046
rect 3045 -5135 3109 -5129
rect 3045 -5251 3051 -5135
rect 3103 -5251 3109 -5135
rect 1513 -5867 1577 -5861
rect 1513 -5983 1519 -5867
rect 1571 -5983 1577 -5867
rect 1513 -6053 1577 -5983
rect 593 -6201 657 -6197
rect 593 -6257 597 -6201
rect 653 -6257 657 -6201
rect 593 -7367 657 -6257
rect 1085 -6270 1149 -6261
rect 1140 -6357 1196 -6352
rect 3045 -6357 3109 -5251
rect 1136 -6361 1200 -6357
rect 1136 -6417 1140 -6361
rect 1196 -6417 1200 -6361
rect 1136 -7332 1200 -6417
rect 3045 -6430 3109 -6421
rect 1669 -6511 1725 -6506
rect 3183 -6511 3247 -5042
rect 5157 -5135 5221 -5129
rect 5157 -5251 5163 -5135
rect 5215 -5251 5221 -5135
rect 3625 -5867 3689 -5861
rect 3625 -5983 3631 -5867
rect 3683 -5983 3689 -5867
rect 3625 -6053 3689 -5983
rect 1665 -6515 1729 -6511
rect 1665 -6571 1669 -6515
rect 1725 -6571 1729 -6515
rect 1665 -7375 1729 -6571
rect 3183 -6584 3247 -6575
rect 2205 -6658 2261 -6653
rect 5157 -6658 5221 -5251
rect 2201 -6662 2265 -6658
rect 2201 -6718 2205 -6662
rect 2261 -6718 2265 -6662
rect 2201 -7382 2265 -6718
rect 5157 -6731 5221 -6722
rect 2747 -6812 2803 -6807
rect 5303 -6812 5367 -5035
rect 7269 -5135 7333 -5129
rect 7269 -5251 7275 -5135
rect 7327 -5251 7333 -5135
rect 5737 -5867 5801 -5861
rect 5737 -5983 5743 -5867
rect 5795 -5983 5801 -5867
rect 5737 -6053 5801 -5983
rect 2743 -6816 2807 -6812
rect 2743 -6872 2747 -6816
rect 2803 -6872 2807 -6816
rect 2743 -7390 2807 -6872
rect 5303 -6885 5367 -6876
rect 3275 -6996 3331 -6991
rect 7269 -6996 7333 -5251
rect 3271 -7000 3335 -6996
rect 3271 -7056 3275 -7000
rect 3331 -7056 3335 -7000
rect 3271 -7368 3335 -7056
rect 7269 -7069 7333 -7060
rect 3805 -7143 3861 -7138
rect 7416 -7143 7480 -5006
rect 9381 -5135 9445 -5129
rect 9381 -5251 9387 -5135
rect 9439 -5251 9445 -5135
rect 7849 -5867 7913 -5861
rect 7849 -5983 7855 -5867
rect 7907 -5983 7913 -5867
rect 7849 -6053 7913 -5983
rect 3801 -7147 3865 -7143
rect 3801 -7203 3805 -7147
rect 3861 -7203 3865 -7147
rect 3801 -7368 3865 -7203
rect 7407 -7207 7416 -7143
rect 7480 -7207 7489 -7143
rect 3961 -7390 4025 -7248
rect -4580 -7700 -4574 -7564
rect -4386 -7700 -4380 -7564
rect 9381 -7520 9445 -5251
rect 9381 -7593 9445 -7584
rect -4580 -7706 -4380 -7700
rect -4390 -8042 -4330 -8033
rect -4390 -8904 -4330 -8102
rect -4390 -8960 -4388 -8904
rect -4332 -8960 -4330 -8904
rect -4390 -8962 -4330 -8960
rect -4388 -8969 -4332 -8962
rect -27806 -10796 -27800 -10519
rect -27412 -10796 -27406 -10519
rect -27806 -10802 -27406 -10796
rect -28262 -11096 -28256 -10858
rect -27868 -11096 -27862 -10858
rect -5082 -10830 -4381 -10824
rect -5082 -11018 -5076 -10830
rect -4893 -11018 -4575 -10830
rect -4387 -11018 -4381 -10830
rect -5082 -11024 -4381 -11018
rect -28262 -11102 -27862 -11096
<< via2 >>
rect -27929 10119 -27868 10255
rect -19249 7687 -19185 7751
rect -27035 7091 -26979 7147
rect -27478 6676 -27412 6812
rect -27478 2178 -27412 2314
rect -17661 7087 -17597 7151
rect -18588 5454 -18528 5514
rect -18293 5250 -18229 5314
rect -4649 1414 -4519 1416
rect -4649 1288 -4647 1414
rect -4647 1288 -4521 1414
rect -4521 1288 -4519 1414
rect -4649 1286 -4519 1288
rect -4435 1340 -4379 1342
rect -4435 1288 -4433 1340
rect -4433 1288 -4381 1340
rect -4381 1288 -4379 1340
rect -4435 1286 -4379 1288
rect -4300 1414 -4244 1416
rect -4300 1288 -4298 1414
rect -4298 1288 -4246 1414
rect -4246 1288 -4244 1414
rect -4300 1286 -4244 1288
rect -5133 1038 -5003 1168
rect -4918 1038 -4862 1094
rect -4784 1038 -4728 1168
rect -4649 1166 -4519 1168
rect -4649 1040 -4647 1166
rect -4647 1040 -4521 1166
rect -4521 1040 -4519 1166
rect -4649 1038 -4519 1040
rect -4435 1092 -4379 1094
rect -4435 1040 -4433 1092
rect -4433 1040 -4381 1092
rect -4381 1040 -4379 1092
rect -4435 1038 -4379 1040
rect -4300 1166 -4244 1168
rect -4300 1040 -4298 1166
rect -4298 1040 -4246 1166
rect -4246 1040 -4244 1166
rect -4300 1038 -4244 1040
rect -4775 758 -4645 814
rect -4291 768 -4161 770
rect -4291 716 -4289 768
rect -4289 716 -4163 768
rect -4163 716 -4161 768
rect -4291 714 -4161 716
rect -12959 -967 -12895 -903
rect -17657 -2734 -17601 -2678
rect -12955 -3434 -12899 -3378
rect -9597 -3438 -9533 -3374
rect -9593 -3746 -9537 -3690
rect -5287 -6940 -5223 -6876
rect -5403 -7078 -5339 -7014
rect -7405 -7216 -7341 -7152
rect -7515 -7362 -7451 -7298
rect -13158 -7580 -13102 -7524
rect -5084 -7580 -5028 -7524
rect -18586 -8100 -18530 -8044
rect -3175 -6608 -3111 -6544
rect -1529 -6604 -1473 -6548
rect -3291 -6774 -3227 -6710
rect -2079 -6770 -2023 -6714
rect -2614 -6936 -2558 -6880
rect -3142 -7074 -3086 -7018
rect -3666 -7212 -3610 -7156
rect -4212 -7358 -4156 -7302
rect 9381 -3750 9445 -3686
rect 76 -6119 132 -6063
rect -1020 -7186 -956 -7122
rect -466 -7182 -410 -7126
rect 933 -6123 997 -6059
rect 597 -6257 653 -6201
rect 1085 -6261 1149 -6197
rect 1140 -6417 1196 -6361
rect 3045 -6421 3109 -6357
rect 1669 -6571 1725 -6515
rect 3183 -6575 3247 -6511
rect 2205 -6718 2261 -6662
rect 5157 -6722 5221 -6658
rect 2747 -6872 2803 -6816
rect 5303 -6876 5367 -6812
rect 3275 -7056 3331 -7000
rect 7269 -7060 7333 -6996
rect 3805 -7203 3861 -7147
rect 7416 -7207 7480 -7143
rect 9381 -7584 9445 -7520
rect -4390 -8102 -4330 -8042
rect -4388 -8960 -4332 -8904
<< metal3 >>
rect -27935 10255 -27136 10261
rect -27935 10119 -27929 10255
rect -27868 10119 -27136 10255
rect -27935 10113 -27136 10119
rect -27218 7751 -19180 7756
rect -27218 7687 -19249 7751
rect -19185 7687 -19180 7751
rect -27218 7682 -19180 7687
rect -27040 7151 -26974 7152
rect -17666 7151 -17592 7156
rect -27040 7147 -17661 7151
rect -27040 7091 -27035 7147
rect -26979 7091 -17661 7147
rect -27040 7087 -17661 7091
rect -17597 7087 -17592 7151
rect -27040 7086 -26974 7087
rect -17666 7082 -17592 7087
rect -27484 6812 -27166 6818
rect -27484 6676 -27478 6812
rect -27412 6676 -27166 6812
rect -27484 6670 -27166 6676
rect -18593 5514 -18523 5519
rect -18593 5454 -18588 5514
rect -18528 5454 -18523 5514
rect -18593 5449 -18523 5454
rect -18298 5314 -18224 5319
rect -18298 5250 -18293 5314
rect -18229 5250 -18224 5314
rect -18298 5245 -18224 5250
rect -27484 2314 -26420 2320
rect -27484 2178 -27478 2314
rect -27412 2178 -26420 2314
rect -27484 2172 -26420 2178
rect -4658 1416 -4510 1425
rect -4658 1286 -4649 1416
rect -4519 1286 -4510 1416
rect -4309 1416 -4235 1425
rect -4658 1277 -4510 1286
rect -4444 1342 -4370 1351
rect -4444 1286 -4435 1342
rect -4379 1286 -4370 1342
rect -4444 1277 -4370 1286
rect -4309 1286 -4300 1416
rect -4244 1286 -4235 1416
rect -4309 1277 -4235 1286
rect -5142 1168 -4994 1177
rect -5142 1038 -5133 1168
rect -5003 1038 -4994 1168
rect -4793 1168 -4719 1177
rect -5142 1029 -4994 1038
rect -4927 1094 -4853 1103
rect -4927 1038 -4918 1094
rect -4862 1038 -4853 1094
rect -4927 1029 -4853 1038
rect -4793 1038 -4784 1168
rect -4728 1038 -4719 1168
rect -4793 1029 -4719 1038
rect -4658 1168 -4510 1177
rect -4658 1038 -4649 1168
rect -4519 1038 -4510 1168
rect -4309 1168 -4235 1177
rect -4658 1029 -4510 1038
rect -4444 1094 -4370 1103
rect -4444 1038 -4435 1094
rect -4379 1038 -4370 1094
rect -4444 1029 -4370 1038
rect -4309 1038 -4300 1168
rect -4244 1038 -4235 1168
rect -4309 1029 -4235 1038
rect -4784 814 -4636 823
rect -4784 758 -4775 814
rect -4645 758 -4636 814
rect -4784 749 -4636 758
rect -4300 770 -4152 779
rect -4300 714 -4291 770
rect -4161 714 -4152 770
rect -4300 705 -4152 714
rect -12964 -903 -12890 -898
rect -12964 -967 -12959 -903
rect -12895 -967 -12890 -903
rect -12964 -972 -12890 -967
rect -17662 -2674 -17596 -2673
rect -17662 -2678 -15348 -2674
rect -17662 -2734 -17657 -2678
rect -17601 -2734 -15348 -2678
rect -17662 -2738 -15348 -2734
rect -17662 -2739 -17596 -2738
rect -15414 -2793 -15348 -2738
rect -15414 -2858 -15412 -2793
rect -12960 -3374 -12894 -3373
rect -9602 -3374 -9528 -3369
rect -12960 -3378 -9597 -3374
rect -12960 -3434 -12955 -3378
rect -12899 -3434 -9597 -3378
rect -12960 -3438 -9597 -3434
rect -9533 -3438 -9528 -3374
rect -12960 -3439 -12894 -3438
rect -9602 -3443 -9528 -3438
rect -9598 -3686 -9532 -3685
rect 9376 -3686 9450 -3681
rect -9598 -3690 9381 -3686
rect -9598 -3746 -9593 -3690
rect -9537 -3746 9381 -3690
rect -9598 -3750 9381 -3746
rect 9445 -3750 9450 -3686
rect -9598 -3751 -9532 -3750
rect 9376 -3755 9450 -3750
rect 71 -6059 137 -6058
rect 928 -6059 1002 -6054
rect 71 -6063 933 -6059
rect 71 -6119 76 -6063
rect 132 -6119 933 -6063
rect 71 -6123 933 -6119
rect 997 -6123 1002 -6059
rect 71 -6124 137 -6123
rect 928 -6128 1002 -6123
rect 592 -6197 658 -6196
rect 1080 -6197 1154 -6192
rect 592 -6201 1085 -6197
rect 592 -6257 597 -6201
rect 653 -6257 1085 -6201
rect 592 -6261 1085 -6257
rect 1149 -6261 1154 -6197
rect 592 -6262 658 -6261
rect 1080 -6266 1154 -6261
rect 1135 -6357 1201 -6356
rect 3040 -6357 3114 -6352
rect 1135 -6361 3045 -6357
rect 1135 -6417 1140 -6361
rect 1196 -6417 3045 -6361
rect 1135 -6421 3045 -6417
rect 3109 -6421 3114 -6357
rect 1135 -6422 1201 -6421
rect 3040 -6426 3114 -6421
rect 1664 -6511 1730 -6510
rect 3178 -6511 3252 -6506
rect 1664 -6515 3183 -6511
rect -3180 -6544 -3106 -6539
rect -1534 -6544 -1468 -6543
rect -3180 -6608 -3175 -6544
rect -3111 -6548 -1468 -6544
rect -3111 -6604 -1529 -6548
rect -1473 -6604 -1468 -6548
rect 1664 -6571 1669 -6515
rect 1725 -6571 3183 -6515
rect 1664 -6575 3183 -6571
rect 3247 -6575 3252 -6511
rect 1664 -6576 1730 -6575
rect 3178 -6580 3252 -6575
rect -3111 -6608 -1468 -6604
rect -3180 -6613 -3106 -6608
rect -1534 -6609 -1468 -6608
rect 2200 -6658 2266 -6657
rect 5152 -6658 5226 -6653
rect 2200 -6662 5157 -6658
rect -3296 -6710 -3222 -6705
rect -2084 -6710 -2018 -6709
rect -3296 -6774 -3291 -6710
rect -3227 -6714 -2018 -6710
rect -3227 -6770 -2079 -6714
rect -2023 -6770 -2018 -6714
rect 2200 -6718 2205 -6662
rect 2261 -6718 5157 -6662
rect 2200 -6722 5157 -6718
rect 5221 -6722 5226 -6658
rect 2200 -6723 2266 -6722
rect 5152 -6727 5226 -6722
rect -3227 -6774 -2018 -6770
rect -3296 -6779 -3222 -6774
rect -2084 -6775 -2018 -6774
rect 2742 -6812 2808 -6811
rect 5298 -6812 5372 -6807
rect 2742 -6816 5303 -6812
rect -5292 -6876 -5218 -6871
rect 2742 -6872 2747 -6816
rect 2803 -6872 5303 -6816
rect -2619 -6876 -2553 -6875
rect -5292 -6940 -5287 -6876
rect -5223 -6880 -2553 -6876
rect 2742 -6876 5303 -6872
rect 5367 -6876 5372 -6812
rect 2742 -6877 2808 -6876
rect -5223 -6936 -2614 -6880
rect -2558 -6936 -2553 -6880
rect 5298 -6881 5372 -6876
rect -5223 -6940 -2553 -6936
rect -5292 -6945 -5218 -6940
rect -2619 -6941 -2553 -6940
rect 3270 -6996 3336 -6995
rect 7264 -6996 7338 -6991
rect 3270 -7000 7269 -6996
rect -5408 -7014 -5334 -7009
rect -3147 -7014 -3081 -7013
rect -5408 -7078 -5403 -7014
rect -5339 -7018 -3081 -7014
rect -5339 -7074 -3142 -7018
rect -3086 -7074 -3081 -7018
rect 3270 -7056 3275 -7000
rect 3331 -7056 7269 -7000
rect 3270 -7060 7269 -7056
rect 7333 -7060 7338 -6996
rect 3270 -7061 3336 -7060
rect 7264 -7065 7338 -7060
rect -5339 -7078 -3081 -7074
rect -5408 -7083 -5334 -7078
rect -3147 -7079 -3081 -7078
rect -1025 -7122 -951 -7117
rect -471 -7122 -405 -7121
rect -7410 -7152 -7336 -7147
rect -3671 -7152 -3605 -7151
rect -7410 -7216 -7405 -7152
rect -7341 -7156 -3605 -7152
rect -7341 -7212 -3666 -7156
rect -3610 -7212 -3605 -7156
rect -1025 -7186 -1020 -7122
rect -956 -7126 -405 -7122
rect -956 -7182 -466 -7126
rect -410 -7182 -405 -7126
rect -956 -7186 -405 -7182
rect -1025 -7191 -951 -7186
rect -471 -7187 -405 -7186
rect 3800 -7143 3866 -7142
rect 7411 -7143 7485 -7138
rect 3800 -7147 7416 -7143
rect 3800 -7203 3805 -7147
rect 3861 -7203 7416 -7147
rect 3800 -7207 7416 -7203
rect 7480 -7207 7485 -7143
rect 3800 -7208 3866 -7207
rect 7411 -7212 7485 -7207
rect -7341 -7216 -3605 -7212
rect -7410 -7221 -7336 -7216
rect -3671 -7217 -3605 -7216
rect -7520 -7298 -7446 -7293
rect -4217 -7298 -4151 -7297
rect -7520 -7362 -7515 -7298
rect -7451 -7302 -4151 -7298
rect -7451 -7358 -4212 -7302
rect -4156 -7358 -4151 -7302
rect -7451 -7362 -4151 -7358
rect -7520 -7367 -7446 -7362
rect -4217 -7363 -4151 -7362
rect -13163 -7520 -13097 -7519
rect -5089 -7520 -5023 -7519
rect 9376 -7520 9450 -7515
rect -13163 -7524 9381 -7520
rect -13163 -7580 -13158 -7524
rect -13102 -7580 -5084 -7524
rect -5028 -7580 9381 -7524
rect -13163 -7584 9381 -7580
rect 9445 -7584 9450 -7520
rect -13163 -7585 -13097 -7584
rect -5089 -7585 -5023 -7584
rect 9376 -7589 9450 -7584
rect -18591 -8042 -18525 -8039
rect -4395 -8042 -4325 -8037
rect -18591 -8044 -4390 -8042
rect -18591 -8100 -18586 -8044
rect -18530 -8100 -4390 -8044
rect -18591 -8102 -4390 -8100
rect -4330 -8102 -4325 -8042
rect -18591 -8105 -18525 -8102
rect -4395 -8107 -4325 -8102
rect -4393 -8902 -4327 -8899
rect -4393 -8904 -3729 -8902
rect -4393 -8960 -4388 -8904
rect -4332 -8960 -3729 -8904
rect -4393 -8962 -3729 -8960
rect 3724 -8962 3784 -8902
rect -4393 -8965 -4327 -8962
use comparator  comparator_0
timestamp 1712334093
transform 1 0 -26517 0 1 2397
box -811 -518 11035 7864
use ibias_gen  ibias_gen_0
timestamp 1712334093
transform 1 0 -27321 0 1 -10450
box -138 -652 15828 11500
use rstring_mux  rstring_mux_0
timestamp 1712334093
transform 1 0 -16753 0 1 -15968
box -11632 -32 28451 9182
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 8 2112 0 1 1734
timestamp 1707688321
transform 1 0 -9540 0 1 -6297
box -66 -43 2178 1671
<< labels >>
flabel metal2 s -9047 -6053 -9047 -6053 0 FreeSans 1200 0 0 0 otrip_decoded[0]
port 3 nsew
flabel metal2 s -6935 -6053 -6935 -6053 0 FreeSans 1200 0 0 0 otrip_decoded[2]
port 4 nsew
flabel metal2 s -4823 -6053 -4823 -6053 0 FreeSans 1200 0 0 0 otrip_decoded[4]
port 5 nsew
flabel metal2 s -2711 -6053 -2711 -6053 0 FreeSans 1200 0 0 0 otrip_decoded[6]
port 6 nsew
flabel metal2 s -599 -6053 -599 -6053 0 FreeSans 1200 0 0 0 otrip_decoded[8]
port 7 nsew
flabel metal2 s 1513 -6053 1513 -6053 0 FreeSans 1200 0 0 0 otrip_decoded[10]
port 8 nsew
flabel metal2 s 3625 -6053 3625 -6053 0 FreeSans 1200 0 0 0 otrip_decoded[12]
port 9 nsew
flabel metal2 s 5737 -6053 5737 -6053 0 FreeSans 1200 0 0 0 otrip_decoded[14]
port 10 nsew
flabel metal2 s 5737 -4319 5737 -4319 0 FreeSans 1200 0 0 0 otrip_decoded[15]
port 11 nsew
flabel metal2 s 3625 -4319 3625 -4319 0 FreeSans 1200 0 0 0 otrip_decoded[13]
port 12 nsew
flabel metal2 s 1513 -4319 1513 -4319 0 FreeSans 1200 0 0 0 otrip_decoded[11]
port 13 nsew
flabel metal2 s -599 -4319 -599 -4319 0 FreeSans 1200 0 0 0 otrip_decoded[9]
port 14 nsew
flabel metal2 s -2711 -4319 -2711 -4319 0 FreeSans 1200 0 0 0 otrip_decoded[7]
port 15 nsew
flabel metal2 s -4823 -4319 -4823 -4319 0 FreeSans 1200 0 0 0 otrip_decoded[5]
port 16 nsew
flabel metal2 s -6935 -4319 -6935 -4319 0 FreeSans 1200 0 0 0 otrip_decoded[3]
port 17 nsew
flabel metal2 s -9047 -4319 -9047 -4319 0 FreeSans 1200 0 0 0 otrip_decoded[1]
port 18 nsew
flabel metal1 s -4836 -6846 -4836 -6846 0 FreeSans 1200 0 0 0 avdd
port 19 nsew
flabel metal1 s -4580 -7558 -4580 -7558 0 FreeSans 1200 0 0 0 avss
port 20 nsew
flabel metal1 s -4836 -6636 -4836 -6636 0 FreeSans 1200 0 0 0 dvdd
port 21 nsew
flabel metal2 s 7849 -6053 7909 -5993 0 FreeSans 1200 0 0 0 ena
port 23 nsew
flabel metal2 s 7849 -4319 7909 -4259 0 FreeSans 1200 0 0 0 isrc_sel
port 24 nsew
flabel metal2 -17531 753 -17531 753 0 FreeSans 1200 0 0 0 itest
port 25 nsew
flabel metal2 s -18241 -2814 -18241 -2814 0 FreeSans 1200 0 0 0 vbg_1v2
port 26 nsew
flabel metal2 -15287 -2068 -15287 -2068 0 FreeSans 1200 0 0 0 ibg_200n
port 27 nsew
flabel metal3 s 3724 -8962 3784 -8902 0 FreeSans 1200 0 0 0 vin
port 22 nsew
<< end >>
