VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__lsbufhv2lv_1
  CLASS BLOCK ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2lv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 8.140 ;
  PIN A
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.630 4.870 1.300 5.200 ;
    END
  END A
  PIN LVPWR
    ANTENNADIFFAREA 1.176500 ;
    PORT
      LAYER nwell ;
        RECT 3.530 1.925 5.000 5.575 ;
      LAYER li1 ;
        RECT 4.130 4.085 4.400 5.415 ;
        RECT 3.780 3.415 4.750 4.085 ;
        RECT 4.130 3.075 4.750 3.415 ;
        RECT 4.130 2.085 4.400 3.075 ;
      LAYER mcon ;
        RECT 4.160 3.105 4.330 3.275 ;
        RECT 4.520 3.105 4.690 3.275 ;
      LAYER met1 ;
        RECT 0.070 3.020 8.090 3.305 ;
    END
  END LVPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.895 6.745 1.485 7.745 ;
        RECT 2.530 5.615 3.120 7.745 ;
      LAYER mcon ;
        RECT 0.925 7.545 1.095 7.715 ;
        RECT 1.285 7.545 1.455 7.715 ;
        RECT 2.560 7.545 2.730 7.715 ;
        RECT 2.920 7.545 3.090 7.715 ;
      LAYER met1 ;
        RECT 0.000 7.515 8.160 7.885 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.895 0.395 1.485 1.395 ;
        RECT 2.570 0.395 3.160 3.910 ;
        RECT 4.130 0.395 4.720 1.515 ;
      LAYER mcon ;
        RECT 0.925 0.425 1.095 0.595 ;
        RECT 1.285 0.425 1.455 0.595 ;
        RECT 2.600 0.425 2.770 0.595 ;
        RECT 2.960 0.425 3.130 0.595 ;
        RECT 4.160 0.425 4.330 0.595 ;
        RECT 4.520 0.425 4.690 0.595 ;
      LAYER met1 ;
        RECT 0.000 0.255 8.160 0.625 ;
    END
  END VGND
  PIN VNB
    ANTENNADIFFAREA 1.387200 ;
    PORT
      LAYER pwell ;
        RECT 1.830 1.625 3.120 4.055 ;
        RECT 1.830 1.585 4.520 1.625 ;
        RECT 0.020 0.215 4.520 1.585 ;
        RECT -0.130 -0.215 8.290 0.215 ;
      LAYER li1 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.115 8.160 0.115 ;
    END
    PORT
      LAYER pwell ;
        RECT -0.130 7.925 8.290 8.355 ;
        RECT 0.020 6.555 3.900 7.925 ;
        RECT 1.830 5.505 3.120 6.555 ;
      LAYER li1 ;
        RECT 0.000 8.055 8.160 8.225 ;
      LAYER mcon ;
        RECT 0.155 8.055 0.325 8.225 ;
        RECT 0.635 8.055 0.805 8.225 ;
        RECT 1.115 8.055 1.285 8.225 ;
        RECT 1.595 8.055 1.765 8.225 ;
        RECT 2.075 8.055 2.245 8.225 ;
        RECT 2.555 8.055 2.725 8.225 ;
        RECT 3.035 8.055 3.205 8.225 ;
        RECT 3.515 8.055 3.685 8.225 ;
        RECT 3.995 8.055 4.165 8.225 ;
        RECT 4.475 8.055 4.645 8.225 ;
        RECT 4.955 8.055 5.125 8.225 ;
        RECT 5.435 8.055 5.605 8.225 ;
        RECT 5.915 8.055 6.085 8.225 ;
        RECT 6.395 8.055 6.565 8.225 ;
        RECT 6.875 8.055 7.045 8.225 ;
        RECT 7.355 8.055 7.525 8.225 ;
        RECT 7.835 8.055 8.005 8.225 ;
      LAYER met1 ;
        RECT 0.000 8.025 8.160 8.255 ;
    END
  END VNB
  PIN VPB
    ANTENNADIFFAREA 0.345100 ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 1.530 6.255 ;
        RECT 7.000 1.885 8.490 6.255 ;
      LAYER li1 ;
        RECT 0.000 3.985 0.885 4.155 ;
        RECT 7.275 3.985 8.160 4.155 ;
      LAYER mcon ;
        RECT 0.155 3.985 0.325 4.155 ;
        RECT 0.635 3.985 0.805 4.155 ;
        RECT 7.355 3.985 7.525 4.155 ;
        RECT 7.835 3.985 8.005 4.155 ;
      LAYER met1 ;
        RECT 0.000 3.955 8.160 4.185 ;
    END
  END VPB
  PIN VPWR
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.130 3.445 0.720 3.675 ;
        RECT 0.130 2.260 0.460 3.445 ;
      LAYER mcon ;
        RECT 0.160 3.475 0.330 3.645 ;
        RECT 0.520 3.475 0.690 3.645 ;
      LAYER met1 ;
        RECT 0.000 3.445 8.160 3.815 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.130 4.695 0.460 5.880 ;
        RECT 0.130 4.465 0.720 4.695 ;
      LAYER mcon ;
        RECT 0.160 4.495 0.330 4.665 ;
        RECT 0.520 4.495 0.690 4.665 ;
      LAYER met1 ;
        RECT 0.000 4.325 8.160 4.695 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER li1 ;
        RECT 3.485 0.735 3.960 3.245 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.170 6.575 0.420 7.060 ;
        RECT 0.170 6.220 1.750 6.575 ;
        RECT 0.950 5.550 1.750 6.220 ;
        RECT 1.470 3.085 1.750 5.550 ;
        RECT 1.920 5.445 2.250 7.455 ;
        RECT 3.480 5.845 3.810 7.455 ;
        RECT 3.290 5.595 5.170 5.845 ;
        RECT 3.290 5.445 3.540 5.595 ;
        RECT 1.920 5.195 3.540 5.445 ;
        RECT 3.710 4.595 3.960 5.415 ;
        RECT 0.630 2.835 1.750 3.085 ;
        RECT 1.920 4.255 3.960 4.595 ;
        RECT 0.950 1.895 1.200 2.590 ;
        RECT 1.445 1.895 1.750 2.235 ;
        RECT 0.170 1.565 1.750 1.895 ;
        RECT 0.170 1.080 0.420 1.565 ;
        RECT 1.920 0.685 2.250 4.255 ;
        RECT 4.920 2.905 5.170 5.595 ;
        RECT 4.570 2.655 5.170 2.905 ;
        RECT 4.570 2.085 4.820 2.655 ;
  END
END sky130_fd_sc_hvl__lsbufhv2lv_1
END LIBRARY

