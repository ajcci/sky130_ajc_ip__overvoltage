magic
tech sky130A
magscale 1 2
timestamp 1711767182
<< nwell >>
rect -5203 -1300 5203 1300
<< mvpmos >>
rect -4945 989 -3345 1073
rect -3287 989 -1687 1073
rect -1629 989 -29 1073
rect 29 989 1629 1073
rect 1687 989 3287 1073
rect 3345 989 4945 1073
rect -4945 740 -3345 824
rect -3287 740 -1687 824
rect -1629 740 -29 824
rect 29 740 1629 824
rect 1687 740 3287 824
rect 3345 740 4945 824
rect -4945 491 -3345 575
rect -3287 491 -1687 575
rect -1629 491 -29 575
rect 29 491 1629 575
rect 1687 491 3287 575
rect 3345 491 4945 575
rect -4945 242 -3345 326
rect -3287 242 -1687 326
rect -1629 242 -29 326
rect 29 242 1629 326
rect 1687 242 3287 326
rect 3345 242 4945 326
rect -4945 -7 -3345 77
rect -3287 -7 -1687 77
rect -1629 -7 -29 77
rect 29 -7 1629 77
rect 1687 -7 3287 77
rect 3345 -7 4945 77
rect -4945 -256 -3345 -172
rect -3287 -256 -1687 -172
rect -1629 -256 -29 -172
rect 29 -256 1629 -172
rect 1687 -256 3287 -172
rect 3345 -256 4945 -172
rect -4945 -505 -3345 -421
rect -3287 -505 -1687 -421
rect -1629 -505 -29 -421
rect 29 -505 1629 -421
rect 1687 -505 3287 -421
rect 3345 -505 4945 -421
rect -4945 -754 -3345 -670
rect -3287 -754 -1687 -670
rect -1629 -754 -29 -670
rect 29 -754 1629 -670
rect 1687 -754 3287 -670
rect 3345 -754 4945 -670
rect -4945 -1003 -3345 -919
rect -3287 -1003 -1687 -919
rect -1629 -1003 -29 -919
rect 29 -1003 1629 -919
rect 1687 -1003 3287 -919
rect 3345 -1003 4945 -919
<< mvpdiff >>
rect -5003 1061 -4945 1073
rect -5003 1001 -4991 1061
rect -4957 1001 -4945 1061
rect -5003 989 -4945 1001
rect -3345 1061 -3287 1073
rect -3345 1001 -3333 1061
rect -3299 1001 -3287 1061
rect -3345 989 -3287 1001
rect -1687 1061 -1629 1073
rect -1687 1001 -1675 1061
rect -1641 1001 -1629 1061
rect -1687 989 -1629 1001
rect -29 1061 29 1073
rect -29 1001 -17 1061
rect 17 1001 29 1061
rect -29 989 29 1001
rect 1629 1061 1687 1073
rect 1629 1001 1641 1061
rect 1675 1001 1687 1061
rect 1629 989 1687 1001
rect 3287 1061 3345 1073
rect 3287 1001 3299 1061
rect 3333 1001 3345 1061
rect 3287 989 3345 1001
rect 4945 1061 5003 1073
rect 4945 1001 4957 1061
rect 4991 1001 5003 1061
rect 4945 989 5003 1001
rect -5003 812 -4945 824
rect -5003 752 -4991 812
rect -4957 752 -4945 812
rect -5003 740 -4945 752
rect -3345 812 -3287 824
rect -3345 752 -3333 812
rect -3299 752 -3287 812
rect -3345 740 -3287 752
rect -1687 812 -1629 824
rect -1687 752 -1675 812
rect -1641 752 -1629 812
rect -1687 740 -1629 752
rect -29 812 29 824
rect -29 752 -17 812
rect 17 752 29 812
rect -29 740 29 752
rect 1629 812 1687 824
rect 1629 752 1641 812
rect 1675 752 1687 812
rect 1629 740 1687 752
rect 3287 812 3345 824
rect 3287 752 3299 812
rect 3333 752 3345 812
rect 3287 740 3345 752
rect 4945 812 5003 824
rect 4945 752 4957 812
rect 4991 752 5003 812
rect 4945 740 5003 752
rect -5003 563 -4945 575
rect -5003 503 -4991 563
rect -4957 503 -4945 563
rect -5003 491 -4945 503
rect -3345 563 -3287 575
rect -3345 503 -3333 563
rect -3299 503 -3287 563
rect -3345 491 -3287 503
rect -1687 563 -1629 575
rect -1687 503 -1675 563
rect -1641 503 -1629 563
rect -1687 491 -1629 503
rect -29 563 29 575
rect -29 503 -17 563
rect 17 503 29 563
rect -29 491 29 503
rect 1629 563 1687 575
rect 1629 503 1641 563
rect 1675 503 1687 563
rect 1629 491 1687 503
rect 3287 563 3345 575
rect 3287 503 3299 563
rect 3333 503 3345 563
rect 3287 491 3345 503
rect 4945 563 5003 575
rect 4945 503 4957 563
rect 4991 503 5003 563
rect 4945 491 5003 503
rect -5003 314 -4945 326
rect -5003 254 -4991 314
rect -4957 254 -4945 314
rect -5003 242 -4945 254
rect -3345 314 -3287 326
rect -3345 254 -3333 314
rect -3299 254 -3287 314
rect -3345 242 -3287 254
rect -1687 314 -1629 326
rect -1687 254 -1675 314
rect -1641 254 -1629 314
rect -1687 242 -1629 254
rect -29 314 29 326
rect -29 254 -17 314
rect 17 254 29 314
rect -29 242 29 254
rect 1629 314 1687 326
rect 1629 254 1641 314
rect 1675 254 1687 314
rect 1629 242 1687 254
rect 3287 314 3345 326
rect 3287 254 3299 314
rect 3333 254 3345 314
rect 3287 242 3345 254
rect 4945 314 5003 326
rect 4945 254 4957 314
rect 4991 254 5003 314
rect 4945 242 5003 254
rect -5003 65 -4945 77
rect -5003 5 -4991 65
rect -4957 5 -4945 65
rect -5003 -7 -4945 5
rect -3345 65 -3287 77
rect -3345 5 -3333 65
rect -3299 5 -3287 65
rect -3345 -7 -3287 5
rect -1687 65 -1629 77
rect -1687 5 -1675 65
rect -1641 5 -1629 65
rect -1687 -7 -1629 5
rect -29 65 29 77
rect -29 5 -17 65
rect 17 5 29 65
rect -29 -7 29 5
rect 1629 65 1687 77
rect 1629 5 1641 65
rect 1675 5 1687 65
rect 1629 -7 1687 5
rect 3287 65 3345 77
rect 3287 5 3299 65
rect 3333 5 3345 65
rect 3287 -7 3345 5
rect 4945 65 5003 77
rect 4945 5 4957 65
rect 4991 5 5003 65
rect 4945 -7 5003 5
rect -5003 -184 -4945 -172
rect -5003 -244 -4991 -184
rect -4957 -244 -4945 -184
rect -5003 -256 -4945 -244
rect -3345 -184 -3287 -172
rect -3345 -244 -3333 -184
rect -3299 -244 -3287 -184
rect -3345 -256 -3287 -244
rect -1687 -184 -1629 -172
rect -1687 -244 -1675 -184
rect -1641 -244 -1629 -184
rect -1687 -256 -1629 -244
rect -29 -184 29 -172
rect -29 -244 -17 -184
rect 17 -244 29 -184
rect -29 -256 29 -244
rect 1629 -184 1687 -172
rect 1629 -244 1641 -184
rect 1675 -244 1687 -184
rect 1629 -256 1687 -244
rect 3287 -184 3345 -172
rect 3287 -244 3299 -184
rect 3333 -244 3345 -184
rect 3287 -256 3345 -244
rect 4945 -184 5003 -172
rect 4945 -244 4957 -184
rect 4991 -244 5003 -184
rect 4945 -256 5003 -244
rect -5003 -433 -4945 -421
rect -5003 -493 -4991 -433
rect -4957 -493 -4945 -433
rect -5003 -505 -4945 -493
rect -3345 -433 -3287 -421
rect -3345 -493 -3333 -433
rect -3299 -493 -3287 -433
rect -3345 -505 -3287 -493
rect -1687 -433 -1629 -421
rect -1687 -493 -1675 -433
rect -1641 -493 -1629 -433
rect -1687 -505 -1629 -493
rect -29 -433 29 -421
rect -29 -493 -17 -433
rect 17 -493 29 -433
rect -29 -505 29 -493
rect 1629 -433 1687 -421
rect 1629 -493 1641 -433
rect 1675 -493 1687 -433
rect 1629 -505 1687 -493
rect 3287 -433 3345 -421
rect 3287 -493 3299 -433
rect 3333 -493 3345 -433
rect 3287 -505 3345 -493
rect 4945 -433 5003 -421
rect 4945 -493 4957 -433
rect 4991 -493 5003 -433
rect 4945 -505 5003 -493
rect -5003 -682 -4945 -670
rect -5003 -742 -4991 -682
rect -4957 -742 -4945 -682
rect -5003 -754 -4945 -742
rect -3345 -682 -3287 -670
rect -3345 -742 -3333 -682
rect -3299 -742 -3287 -682
rect -3345 -754 -3287 -742
rect -1687 -682 -1629 -670
rect -1687 -742 -1675 -682
rect -1641 -742 -1629 -682
rect -1687 -754 -1629 -742
rect -29 -682 29 -670
rect -29 -742 -17 -682
rect 17 -742 29 -682
rect -29 -754 29 -742
rect 1629 -682 1687 -670
rect 1629 -742 1641 -682
rect 1675 -742 1687 -682
rect 1629 -754 1687 -742
rect 3287 -682 3345 -670
rect 3287 -742 3299 -682
rect 3333 -742 3345 -682
rect 3287 -754 3345 -742
rect 4945 -682 5003 -670
rect 4945 -742 4957 -682
rect 4991 -742 5003 -682
rect 4945 -754 5003 -742
rect -5003 -931 -4945 -919
rect -5003 -991 -4991 -931
rect -4957 -991 -4945 -931
rect -5003 -1003 -4945 -991
rect -3345 -931 -3287 -919
rect -3345 -991 -3333 -931
rect -3299 -991 -3287 -931
rect -3345 -1003 -3287 -991
rect -1687 -931 -1629 -919
rect -1687 -991 -1675 -931
rect -1641 -991 -1629 -931
rect -1687 -1003 -1629 -991
rect -29 -931 29 -919
rect -29 -991 -17 -931
rect 17 -991 29 -931
rect -29 -1003 29 -991
rect 1629 -931 1687 -919
rect 1629 -991 1641 -931
rect 1675 -991 1687 -931
rect 1629 -1003 1687 -991
rect 3287 -931 3345 -919
rect 3287 -991 3299 -931
rect 3333 -991 3345 -931
rect 3287 -1003 3345 -991
rect 4945 -931 5003 -919
rect 4945 -991 4957 -931
rect 4991 -991 5003 -931
rect 4945 -1003 5003 -991
<< mvpdiffc >>
rect -4991 1001 -4957 1061
rect -3333 1001 -3299 1061
rect -1675 1001 -1641 1061
rect -17 1001 17 1061
rect 1641 1001 1675 1061
rect 3299 1001 3333 1061
rect 4957 1001 4991 1061
rect -4991 752 -4957 812
rect -3333 752 -3299 812
rect -1675 752 -1641 812
rect -17 752 17 812
rect 1641 752 1675 812
rect 3299 752 3333 812
rect 4957 752 4991 812
rect -4991 503 -4957 563
rect -3333 503 -3299 563
rect -1675 503 -1641 563
rect -17 503 17 563
rect 1641 503 1675 563
rect 3299 503 3333 563
rect 4957 503 4991 563
rect -4991 254 -4957 314
rect -3333 254 -3299 314
rect -1675 254 -1641 314
rect -17 254 17 314
rect 1641 254 1675 314
rect 3299 254 3333 314
rect 4957 254 4991 314
rect -4991 5 -4957 65
rect -3333 5 -3299 65
rect -1675 5 -1641 65
rect -17 5 17 65
rect 1641 5 1675 65
rect 3299 5 3333 65
rect 4957 5 4991 65
rect -4991 -244 -4957 -184
rect -3333 -244 -3299 -184
rect -1675 -244 -1641 -184
rect -17 -244 17 -184
rect 1641 -244 1675 -184
rect 3299 -244 3333 -184
rect 4957 -244 4991 -184
rect -4991 -493 -4957 -433
rect -3333 -493 -3299 -433
rect -1675 -493 -1641 -433
rect -17 -493 17 -433
rect 1641 -493 1675 -433
rect 3299 -493 3333 -433
rect 4957 -493 4991 -433
rect -4991 -742 -4957 -682
rect -3333 -742 -3299 -682
rect -1675 -742 -1641 -682
rect -17 -742 17 -682
rect 1641 -742 1675 -682
rect 3299 -742 3333 -682
rect 4957 -742 4991 -682
rect -4991 -991 -4957 -931
rect -3333 -991 -3299 -931
rect -1675 -991 -1641 -931
rect -17 -991 17 -931
rect 1641 -991 1675 -931
rect 3299 -991 3333 -931
rect 4957 -991 4991 -931
<< mvnsubdiff >>
rect -5137 1222 5137 1234
rect -5137 1188 -5029 1222
rect 5029 1188 5137 1222
rect -5137 1176 5137 1188
rect -5137 1126 -5079 1176
rect -5137 -1126 -5125 1126
rect -5091 -1126 -5079 1126
rect 5079 1126 5137 1176
rect -5137 -1176 -5079 -1126
rect 5079 -1126 5091 1126
rect 5125 -1126 5137 1126
rect 5079 -1176 5137 -1126
rect -5137 -1188 5137 -1176
rect -5137 -1222 -5029 -1188
rect 5029 -1222 5137 -1188
rect -5137 -1234 5137 -1222
<< mvnsubdiffcont >>
rect -5029 1188 5029 1222
rect -5125 -1126 -5091 1126
rect 5091 -1126 5125 1126
rect -5029 -1222 5029 -1188
<< poly >>
rect -4945 1073 -3345 1099
rect -3287 1073 -1687 1099
rect -1629 1073 -29 1099
rect 29 1073 1629 1099
rect 1687 1073 3287 1099
rect 3345 1073 4945 1099
rect -4945 942 -3345 989
rect -4945 908 -4929 942
rect -3361 908 -3345 942
rect -4945 892 -3345 908
rect -3287 942 -1687 989
rect -3287 908 -3271 942
rect -1703 908 -1687 942
rect -3287 892 -1687 908
rect -1629 942 -29 989
rect -1629 908 -1613 942
rect -45 908 -29 942
rect -1629 892 -29 908
rect 29 942 1629 989
rect 29 908 45 942
rect 1613 908 1629 942
rect 29 892 1629 908
rect 1687 942 3287 989
rect 1687 908 1703 942
rect 3271 908 3287 942
rect 1687 892 3287 908
rect 3345 942 4945 989
rect 3345 908 3361 942
rect 4929 908 4945 942
rect 3345 892 4945 908
rect -4945 824 -3345 850
rect -3287 824 -1687 850
rect -1629 824 -29 850
rect 29 824 1629 850
rect 1687 824 3287 850
rect 3345 824 4945 850
rect -4945 693 -3345 740
rect -4945 659 -4929 693
rect -3361 659 -3345 693
rect -4945 643 -3345 659
rect -3287 693 -1687 740
rect -3287 659 -3271 693
rect -1703 659 -1687 693
rect -3287 643 -1687 659
rect -1629 693 -29 740
rect -1629 659 -1613 693
rect -45 659 -29 693
rect -1629 643 -29 659
rect 29 693 1629 740
rect 29 659 45 693
rect 1613 659 1629 693
rect 29 643 1629 659
rect 1687 693 3287 740
rect 1687 659 1703 693
rect 3271 659 3287 693
rect 1687 643 3287 659
rect 3345 693 4945 740
rect 3345 659 3361 693
rect 4929 659 4945 693
rect 3345 643 4945 659
rect -4945 575 -3345 601
rect -3287 575 -1687 601
rect -1629 575 -29 601
rect 29 575 1629 601
rect 1687 575 3287 601
rect 3345 575 4945 601
rect -4945 444 -3345 491
rect -4945 410 -4929 444
rect -3361 410 -3345 444
rect -4945 394 -3345 410
rect -3287 444 -1687 491
rect -3287 410 -3271 444
rect -1703 410 -1687 444
rect -3287 394 -1687 410
rect -1629 444 -29 491
rect -1629 410 -1613 444
rect -45 410 -29 444
rect -1629 394 -29 410
rect 29 444 1629 491
rect 29 410 45 444
rect 1613 410 1629 444
rect 29 394 1629 410
rect 1687 444 3287 491
rect 1687 410 1703 444
rect 3271 410 3287 444
rect 1687 394 3287 410
rect 3345 444 4945 491
rect 3345 410 3361 444
rect 4929 410 4945 444
rect 3345 394 4945 410
rect -4945 326 -3345 352
rect -3287 326 -1687 352
rect -1629 326 -29 352
rect 29 326 1629 352
rect 1687 326 3287 352
rect 3345 326 4945 352
rect -4945 195 -3345 242
rect -4945 161 -4929 195
rect -3361 161 -3345 195
rect -4945 145 -3345 161
rect -3287 195 -1687 242
rect -3287 161 -3271 195
rect -1703 161 -1687 195
rect -3287 145 -1687 161
rect -1629 195 -29 242
rect -1629 161 -1613 195
rect -45 161 -29 195
rect -1629 145 -29 161
rect 29 195 1629 242
rect 29 161 45 195
rect 1613 161 1629 195
rect 29 145 1629 161
rect 1687 195 3287 242
rect 1687 161 1703 195
rect 3271 161 3287 195
rect 1687 145 3287 161
rect 3345 195 4945 242
rect 3345 161 3361 195
rect 4929 161 4945 195
rect 3345 145 4945 161
rect -4945 77 -3345 103
rect -3287 77 -1687 103
rect -1629 77 -29 103
rect 29 77 1629 103
rect 1687 77 3287 103
rect 3345 77 4945 103
rect -4945 -54 -3345 -7
rect -4945 -88 -4929 -54
rect -3361 -88 -3345 -54
rect -4945 -104 -3345 -88
rect -3287 -54 -1687 -7
rect -3287 -88 -3271 -54
rect -1703 -88 -1687 -54
rect -3287 -104 -1687 -88
rect -1629 -54 -29 -7
rect -1629 -88 -1613 -54
rect -45 -88 -29 -54
rect -1629 -104 -29 -88
rect 29 -54 1629 -7
rect 29 -88 45 -54
rect 1613 -88 1629 -54
rect 29 -104 1629 -88
rect 1687 -54 3287 -7
rect 1687 -88 1703 -54
rect 3271 -88 3287 -54
rect 1687 -104 3287 -88
rect 3345 -54 4945 -7
rect 3345 -88 3361 -54
rect 4929 -88 4945 -54
rect 3345 -104 4945 -88
rect -4945 -172 -3345 -146
rect -3287 -172 -1687 -146
rect -1629 -172 -29 -146
rect 29 -172 1629 -146
rect 1687 -172 3287 -146
rect 3345 -172 4945 -146
rect -4945 -303 -3345 -256
rect -4945 -337 -4929 -303
rect -3361 -337 -3345 -303
rect -4945 -353 -3345 -337
rect -3287 -303 -1687 -256
rect -3287 -337 -3271 -303
rect -1703 -337 -1687 -303
rect -3287 -353 -1687 -337
rect -1629 -303 -29 -256
rect -1629 -337 -1613 -303
rect -45 -337 -29 -303
rect -1629 -353 -29 -337
rect 29 -303 1629 -256
rect 29 -337 45 -303
rect 1613 -337 1629 -303
rect 29 -353 1629 -337
rect 1687 -303 3287 -256
rect 1687 -337 1703 -303
rect 3271 -337 3287 -303
rect 1687 -353 3287 -337
rect 3345 -303 4945 -256
rect 3345 -337 3361 -303
rect 4929 -337 4945 -303
rect 3345 -353 4945 -337
rect -4945 -421 -3345 -395
rect -3287 -421 -1687 -395
rect -1629 -421 -29 -395
rect 29 -421 1629 -395
rect 1687 -421 3287 -395
rect 3345 -421 4945 -395
rect -4945 -552 -3345 -505
rect -4945 -586 -4929 -552
rect -3361 -586 -3345 -552
rect -4945 -602 -3345 -586
rect -3287 -552 -1687 -505
rect -3287 -586 -3271 -552
rect -1703 -586 -1687 -552
rect -3287 -602 -1687 -586
rect -1629 -552 -29 -505
rect -1629 -586 -1613 -552
rect -45 -586 -29 -552
rect -1629 -602 -29 -586
rect 29 -552 1629 -505
rect 29 -586 45 -552
rect 1613 -586 1629 -552
rect 29 -602 1629 -586
rect 1687 -552 3287 -505
rect 1687 -586 1703 -552
rect 3271 -586 3287 -552
rect 1687 -602 3287 -586
rect 3345 -552 4945 -505
rect 3345 -586 3361 -552
rect 4929 -586 4945 -552
rect 3345 -602 4945 -586
rect -4945 -670 -3345 -644
rect -3287 -670 -1687 -644
rect -1629 -670 -29 -644
rect 29 -670 1629 -644
rect 1687 -670 3287 -644
rect 3345 -670 4945 -644
rect -4945 -801 -3345 -754
rect -4945 -835 -4929 -801
rect -3361 -835 -3345 -801
rect -4945 -851 -3345 -835
rect -3287 -801 -1687 -754
rect -3287 -835 -3271 -801
rect -1703 -835 -1687 -801
rect -3287 -851 -1687 -835
rect -1629 -801 -29 -754
rect -1629 -835 -1613 -801
rect -45 -835 -29 -801
rect -1629 -851 -29 -835
rect 29 -801 1629 -754
rect 29 -835 45 -801
rect 1613 -835 1629 -801
rect 29 -851 1629 -835
rect 1687 -801 3287 -754
rect 1687 -835 1703 -801
rect 3271 -835 3287 -801
rect 1687 -851 3287 -835
rect 3345 -801 4945 -754
rect 3345 -835 3361 -801
rect 4929 -835 4945 -801
rect 3345 -851 4945 -835
rect -4945 -919 -3345 -893
rect -3287 -919 -1687 -893
rect -1629 -919 -29 -893
rect 29 -919 1629 -893
rect 1687 -919 3287 -893
rect 3345 -919 4945 -893
rect -4945 -1050 -3345 -1003
rect -4945 -1084 -4929 -1050
rect -3361 -1084 -3345 -1050
rect -4945 -1100 -3345 -1084
rect -3287 -1050 -1687 -1003
rect -3287 -1084 -3271 -1050
rect -1703 -1084 -1687 -1050
rect -3287 -1100 -1687 -1084
rect -1629 -1050 -29 -1003
rect -1629 -1084 -1613 -1050
rect -45 -1084 -29 -1050
rect -1629 -1100 -29 -1084
rect 29 -1050 1629 -1003
rect 29 -1084 45 -1050
rect 1613 -1084 1629 -1050
rect 29 -1100 1629 -1084
rect 1687 -1050 3287 -1003
rect 1687 -1084 1703 -1050
rect 3271 -1084 3287 -1050
rect 1687 -1100 3287 -1084
rect 3345 -1050 4945 -1003
rect 3345 -1084 3361 -1050
rect 4929 -1084 4945 -1050
rect 3345 -1100 4945 -1084
<< polycont >>
rect -4929 908 -3361 942
rect -3271 908 -1703 942
rect -1613 908 -45 942
rect 45 908 1613 942
rect 1703 908 3271 942
rect 3361 908 4929 942
rect -4929 659 -3361 693
rect -3271 659 -1703 693
rect -1613 659 -45 693
rect 45 659 1613 693
rect 1703 659 3271 693
rect 3361 659 4929 693
rect -4929 410 -3361 444
rect -3271 410 -1703 444
rect -1613 410 -45 444
rect 45 410 1613 444
rect 1703 410 3271 444
rect 3361 410 4929 444
rect -4929 161 -3361 195
rect -3271 161 -1703 195
rect -1613 161 -45 195
rect 45 161 1613 195
rect 1703 161 3271 195
rect 3361 161 4929 195
rect -4929 -88 -3361 -54
rect -3271 -88 -1703 -54
rect -1613 -88 -45 -54
rect 45 -88 1613 -54
rect 1703 -88 3271 -54
rect 3361 -88 4929 -54
rect -4929 -337 -3361 -303
rect -3271 -337 -1703 -303
rect -1613 -337 -45 -303
rect 45 -337 1613 -303
rect 1703 -337 3271 -303
rect 3361 -337 4929 -303
rect -4929 -586 -3361 -552
rect -3271 -586 -1703 -552
rect -1613 -586 -45 -552
rect 45 -586 1613 -552
rect 1703 -586 3271 -552
rect 3361 -586 4929 -552
rect -4929 -835 -3361 -801
rect -3271 -835 -1703 -801
rect -1613 -835 -45 -801
rect 45 -835 1613 -801
rect 1703 -835 3271 -801
rect 3361 -835 4929 -801
rect -4929 -1084 -3361 -1050
rect -3271 -1084 -1703 -1050
rect -1613 -1084 -45 -1050
rect 45 -1084 1613 -1050
rect 1703 -1084 3271 -1050
rect 3361 -1084 4929 -1050
<< locali >>
rect -5125 1188 -5029 1222
rect 5029 1188 5125 1222
rect -5125 1126 -5091 1188
rect 5091 1126 5125 1188
rect -4991 1061 -4957 1077
rect -4991 985 -4957 1001
rect -3333 1061 -3299 1077
rect -3333 985 -3299 1001
rect -1675 1061 -1641 1077
rect -1675 985 -1641 1001
rect -17 1061 17 1077
rect -17 985 17 1001
rect 1641 1061 1675 1077
rect 1641 985 1675 1001
rect 3299 1061 3333 1077
rect 3299 985 3333 1001
rect 4957 1061 4991 1077
rect 4957 985 4991 1001
rect -4945 908 -4929 942
rect -3361 908 -3345 942
rect -3287 908 -3271 942
rect -1703 908 -1687 942
rect -1629 908 -1613 942
rect -45 908 -29 942
rect 29 908 45 942
rect 1613 908 1629 942
rect 1687 908 1703 942
rect 3271 908 3287 942
rect 3345 908 3361 942
rect 4929 908 4945 942
rect -4991 812 -4957 828
rect -4991 736 -4957 752
rect -3333 812 -3299 828
rect -3333 736 -3299 752
rect -1675 812 -1641 828
rect -1675 736 -1641 752
rect -17 812 17 828
rect -17 736 17 752
rect 1641 812 1675 828
rect 1641 736 1675 752
rect 3299 812 3333 828
rect 3299 736 3333 752
rect 4957 812 4991 828
rect 4957 736 4991 752
rect -4945 659 -4929 693
rect -3361 659 -3345 693
rect -3287 659 -3271 693
rect -1703 659 -1687 693
rect -1629 659 -1613 693
rect -45 659 -29 693
rect 29 659 45 693
rect 1613 659 1629 693
rect 1687 659 1703 693
rect 3271 659 3287 693
rect 3345 659 3361 693
rect 4929 659 4945 693
rect -4991 563 -4957 579
rect -4991 487 -4957 503
rect -3333 563 -3299 579
rect -3333 487 -3299 503
rect -1675 563 -1641 579
rect -1675 487 -1641 503
rect -17 563 17 579
rect -17 487 17 503
rect 1641 563 1675 579
rect 1641 487 1675 503
rect 3299 563 3333 579
rect 3299 487 3333 503
rect 4957 563 4991 579
rect 4957 487 4991 503
rect -4945 410 -4929 444
rect -3361 410 -3345 444
rect -3287 410 -3271 444
rect -1703 410 -1687 444
rect -1629 410 -1613 444
rect -45 410 -29 444
rect 29 410 45 444
rect 1613 410 1629 444
rect 1687 410 1703 444
rect 3271 410 3287 444
rect 3345 410 3361 444
rect 4929 410 4945 444
rect -4991 314 -4957 330
rect -4991 238 -4957 254
rect -3333 314 -3299 330
rect -3333 238 -3299 254
rect -1675 314 -1641 330
rect -1675 238 -1641 254
rect -17 314 17 330
rect -17 238 17 254
rect 1641 314 1675 330
rect 1641 238 1675 254
rect 3299 314 3333 330
rect 3299 238 3333 254
rect 4957 314 4991 330
rect 4957 238 4991 254
rect -4945 161 -4929 195
rect -3361 161 -3345 195
rect -3287 161 -3271 195
rect -1703 161 -1687 195
rect -1629 161 -1613 195
rect -45 161 -29 195
rect 29 161 45 195
rect 1613 161 1629 195
rect 1687 161 1703 195
rect 3271 161 3287 195
rect 3345 161 3361 195
rect 4929 161 4945 195
rect -4991 65 -4957 81
rect -4991 -11 -4957 5
rect -3333 65 -3299 81
rect -3333 -11 -3299 5
rect -1675 65 -1641 81
rect -1675 -11 -1641 5
rect -17 65 17 81
rect -17 -11 17 5
rect 1641 65 1675 81
rect 1641 -11 1675 5
rect 3299 65 3333 81
rect 3299 -11 3333 5
rect 4957 65 4991 81
rect 4957 -11 4991 5
rect -4945 -88 -4929 -54
rect -3361 -88 -3345 -54
rect -3287 -88 -3271 -54
rect -1703 -88 -1687 -54
rect -1629 -88 -1613 -54
rect -45 -88 -29 -54
rect 29 -88 45 -54
rect 1613 -88 1629 -54
rect 1687 -88 1703 -54
rect 3271 -88 3287 -54
rect 3345 -88 3361 -54
rect 4929 -88 4945 -54
rect -4991 -184 -4957 -168
rect -4991 -260 -4957 -244
rect -3333 -184 -3299 -168
rect -3333 -260 -3299 -244
rect -1675 -184 -1641 -168
rect -1675 -260 -1641 -244
rect -17 -184 17 -168
rect -17 -260 17 -244
rect 1641 -184 1675 -168
rect 1641 -260 1675 -244
rect 3299 -184 3333 -168
rect 3299 -260 3333 -244
rect 4957 -184 4991 -168
rect 4957 -260 4991 -244
rect -4945 -337 -4929 -303
rect -3361 -337 -3345 -303
rect -3287 -337 -3271 -303
rect -1703 -337 -1687 -303
rect -1629 -337 -1613 -303
rect -45 -337 -29 -303
rect 29 -337 45 -303
rect 1613 -337 1629 -303
rect 1687 -337 1703 -303
rect 3271 -337 3287 -303
rect 3345 -337 3361 -303
rect 4929 -337 4945 -303
rect -4991 -433 -4957 -417
rect -4991 -509 -4957 -493
rect -3333 -433 -3299 -417
rect -3333 -509 -3299 -493
rect -1675 -433 -1641 -417
rect -1675 -509 -1641 -493
rect -17 -433 17 -417
rect -17 -509 17 -493
rect 1641 -433 1675 -417
rect 1641 -509 1675 -493
rect 3299 -433 3333 -417
rect 3299 -509 3333 -493
rect 4957 -433 4991 -417
rect 4957 -509 4991 -493
rect -4945 -586 -4929 -552
rect -3361 -586 -3345 -552
rect -3287 -586 -3271 -552
rect -1703 -586 -1687 -552
rect -1629 -586 -1613 -552
rect -45 -586 -29 -552
rect 29 -586 45 -552
rect 1613 -586 1629 -552
rect 1687 -586 1703 -552
rect 3271 -586 3287 -552
rect 3345 -586 3361 -552
rect 4929 -586 4945 -552
rect -4991 -682 -4957 -666
rect -4991 -758 -4957 -742
rect -3333 -682 -3299 -666
rect -3333 -758 -3299 -742
rect -1675 -682 -1641 -666
rect -1675 -758 -1641 -742
rect -17 -682 17 -666
rect -17 -758 17 -742
rect 1641 -682 1675 -666
rect 1641 -758 1675 -742
rect 3299 -682 3333 -666
rect 3299 -758 3333 -742
rect 4957 -682 4991 -666
rect 4957 -758 4991 -742
rect -4945 -835 -4929 -801
rect -3361 -835 -3345 -801
rect -3287 -835 -3271 -801
rect -1703 -835 -1687 -801
rect -1629 -835 -1613 -801
rect -45 -835 -29 -801
rect 29 -835 45 -801
rect 1613 -835 1629 -801
rect 1687 -835 1703 -801
rect 3271 -835 3287 -801
rect 3345 -835 3361 -801
rect 4929 -835 4945 -801
rect -4991 -931 -4957 -915
rect -4991 -1007 -4957 -991
rect -3333 -931 -3299 -915
rect -3333 -1007 -3299 -991
rect -1675 -931 -1641 -915
rect -1675 -1007 -1641 -991
rect -17 -931 17 -915
rect -17 -1007 17 -991
rect 1641 -931 1675 -915
rect 1641 -1007 1675 -991
rect 3299 -931 3333 -915
rect 3299 -1007 3333 -991
rect 4957 -931 4991 -915
rect 4957 -1007 4991 -991
rect -4945 -1084 -4929 -1050
rect -3361 -1084 -3345 -1050
rect -3287 -1084 -3271 -1050
rect -1703 -1084 -1687 -1050
rect -1629 -1084 -1613 -1050
rect -45 -1084 -29 -1050
rect 29 -1084 45 -1050
rect 1613 -1084 1629 -1050
rect 1687 -1084 1703 -1050
rect 3271 -1084 3287 -1050
rect 3345 -1084 3361 -1050
rect 4929 -1084 4945 -1050
rect -5125 -1188 -5091 -1126
rect 5091 -1188 5125 -1126
rect -5125 -1222 -5029 -1188
rect 5029 -1222 5125 -1188
<< viali >>
rect -4991 1001 -4957 1061
rect -3333 1001 -3299 1061
rect -1675 1001 -1641 1061
rect -17 1001 17 1061
rect 1641 1001 1675 1061
rect 3299 1001 3333 1061
rect 4957 1001 4991 1061
rect -4929 908 -3361 942
rect -3271 908 -1703 942
rect -1613 908 -45 942
rect 45 908 1613 942
rect 1703 908 3271 942
rect 3361 908 4929 942
rect -4991 752 -4957 812
rect -3333 752 -3299 812
rect -1675 752 -1641 812
rect -17 752 17 812
rect 1641 752 1675 812
rect 3299 752 3333 812
rect 4957 752 4991 812
rect -4929 659 -3361 693
rect -3271 659 -1703 693
rect -1613 659 -45 693
rect 45 659 1613 693
rect 1703 659 3271 693
rect 3361 659 4929 693
rect -4991 503 -4957 563
rect -3333 503 -3299 563
rect -1675 503 -1641 563
rect -17 503 17 563
rect 1641 503 1675 563
rect 3299 503 3333 563
rect 4957 503 4991 563
rect -4929 410 -3361 444
rect -3271 410 -1703 444
rect -1613 410 -45 444
rect 45 410 1613 444
rect 1703 410 3271 444
rect 3361 410 4929 444
rect -4991 254 -4957 314
rect -3333 254 -3299 314
rect -1675 254 -1641 314
rect -17 254 17 314
rect 1641 254 1675 314
rect 3299 254 3333 314
rect 4957 254 4991 314
rect -4929 161 -3361 195
rect -3271 161 -1703 195
rect -1613 161 -45 195
rect 45 161 1613 195
rect 1703 161 3271 195
rect 3361 161 4929 195
rect -4991 5 -4957 65
rect -3333 5 -3299 65
rect -1675 5 -1641 65
rect -17 5 17 65
rect 1641 5 1675 65
rect 3299 5 3333 65
rect 4957 5 4991 65
rect -4929 -88 -3361 -54
rect -3271 -88 -1703 -54
rect -1613 -88 -45 -54
rect 45 -88 1613 -54
rect 1703 -88 3271 -54
rect 3361 -88 4929 -54
rect -4991 -244 -4957 -184
rect -3333 -244 -3299 -184
rect -1675 -244 -1641 -184
rect -17 -244 17 -184
rect 1641 -244 1675 -184
rect 3299 -244 3333 -184
rect 4957 -244 4991 -184
rect -4929 -337 -3361 -303
rect -3271 -337 -1703 -303
rect -1613 -337 -45 -303
rect 45 -337 1613 -303
rect 1703 -337 3271 -303
rect 3361 -337 4929 -303
rect -4991 -493 -4957 -433
rect -3333 -493 -3299 -433
rect -1675 -493 -1641 -433
rect -17 -493 17 -433
rect 1641 -493 1675 -433
rect 3299 -493 3333 -433
rect 4957 -493 4991 -433
rect -4929 -586 -3361 -552
rect -3271 -586 -1703 -552
rect -1613 -586 -45 -552
rect 45 -586 1613 -552
rect 1703 -586 3271 -552
rect 3361 -586 4929 -552
rect -4991 -742 -4957 -682
rect -3333 -742 -3299 -682
rect -1675 -742 -1641 -682
rect -17 -742 17 -682
rect 1641 -742 1675 -682
rect 3299 -742 3333 -682
rect 4957 -742 4991 -682
rect -4929 -835 -3361 -801
rect -3271 -835 -1703 -801
rect -1613 -835 -45 -801
rect 45 -835 1613 -801
rect 1703 -835 3271 -801
rect 3361 -835 4929 -801
rect -4991 -991 -4957 -931
rect -3333 -991 -3299 -931
rect -1675 -991 -1641 -931
rect -17 -991 17 -931
rect 1641 -991 1675 -931
rect 3299 -991 3333 -931
rect 4957 -991 4991 -931
rect -4929 -1084 -3361 -1050
rect -3271 -1084 -1703 -1050
rect -1613 -1084 -45 -1050
rect 45 -1084 1613 -1050
rect 1703 -1084 3271 -1050
rect 3361 -1084 4929 -1050
<< metal1 >>
rect -4997 1061 -4951 1073
rect -4997 1001 -4991 1061
rect -4957 1001 -4951 1061
rect -4997 989 -4951 1001
rect -3339 1061 -3293 1073
rect -3339 1001 -3333 1061
rect -3299 1001 -3293 1061
rect -3339 989 -3293 1001
rect -1681 1061 -1635 1073
rect -1681 1001 -1675 1061
rect -1641 1001 -1635 1061
rect -1681 989 -1635 1001
rect -23 1061 23 1073
rect -23 1001 -17 1061
rect 17 1001 23 1061
rect -23 989 23 1001
rect 1635 1061 1681 1073
rect 1635 1001 1641 1061
rect 1675 1001 1681 1061
rect 1635 989 1681 1001
rect 3293 1061 3339 1073
rect 3293 1001 3299 1061
rect 3333 1001 3339 1061
rect 3293 989 3339 1001
rect 4951 1061 4997 1073
rect 4951 1001 4957 1061
rect 4991 1001 4997 1061
rect 4951 989 4997 1001
rect -4941 942 -3349 948
rect -4941 908 -4929 942
rect -3361 908 -3349 942
rect -4941 902 -3349 908
rect -3283 942 -1691 948
rect -3283 908 -3271 942
rect -1703 908 -1691 942
rect -3283 902 -1691 908
rect -1625 942 -33 948
rect -1625 908 -1613 942
rect -45 908 -33 942
rect -1625 902 -33 908
rect 33 942 1625 948
rect 33 908 45 942
rect 1613 908 1625 942
rect 33 902 1625 908
rect 1691 942 3283 948
rect 1691 908 1703 942
rect 3271 908 3283 942
rect 1691 902 3283 908
rect 3349 942 4941 948
rect 3349 908 3361 942
rect 4929 908 4941 942
rect 3349 902 4941 908
rect -4997 812 -4951 824
rect -4997 752 -4991 812
rect -4957 752 -4951 812
rect -4997 740 -4951 752
rect -3339 812 -3293 824
rect -3339 752 -3333 812
rect -3299 752 -3293 812
rect -3339 740 -3293 752
rect -1681 812 -1635 824
rect -1681 752 -1675 812
rect -1641 752 -1635 812
rect -1681 740 -1635 752
rect -23 812 23 824
rect -23 752 -17 812
rect 17 752 23 812
rect -23 740 23 752
rect 1635 812 1681 824
rect 1635 752 1641 812
rect 1675 752 1681 812
rect 1635 740 1681 752
rect 3293 812 3339 824
rect 3293 752 3299 812
rect 3333 752 3339 812
rect 3293 740 3339 752
rect 4951 812 4997 824
rect 4951 752 4957 812
rect 4991 752 4997 812
rect 4951 740 4997 752
rect -4941 693 -3349 699
rect -4941 659 -4929 693
rect -3361 659 -3349 693
rect -4941 653 -3349 659
rect -3283 693 -1691 699
rect -3283 659 -3271 693
rect -1703 659 -1691 693
rect -3283 653 -1691 659
rect -1625 693 -33 699
rect -1625 659 -1613 693
rect -45 659 -33 693
rect -1625 653 -33 659
rect 33 693 1625 699
rect 33 659 45 693
rect 1613 659 1625 693
rect 33 653 1625 659
rect 1691 693 3283 699
rect 1691 659 1703 693
rect 3271 659 3283 693
rect 1691 653 3283 659
rect 3349 693 4941 699
rect 3349 659 3361 693
rect 4929 659 4941 693
rect 3349 653 4941 659
rect -4997 563 -4951 575
rect -4997 503 -4991 563
rect -4957 503 -4951 563
rect -4997 491 -4951 503
rect -3339 563 -3293 575
rect -3339 503 -3333 563
rect -3299 503 -3293 563
rect -3339 491 -3293 503
rect -1681 563 -1635 575
rect -1681 503 -1675 563
rect -1641 503 -1635 563
rect -1681 491 -1635 503
rect -23 563 23 575
rect -23 503 -17 563
rect 17 503 23 563
rect -23 491 23 503
rect 1635 563 1681 575
rect 1635 503 1641 563
rect 1675 503 1681 563
rect 1635 491 1681 503
rect 3293 563 3339 575
rect 3293 503 3299 563
rect 3333 503 3339 563
rect 3293 491 3339 503
rect 4951 563 4997 575
rect 4951 503 4957 563
rect 4991 503 4997 563
rect 4951 491 4997 503
rect -4941 444 -3349 450
rect -4941 410 -4929 444
rect -3361 410 -3349 444
rect -4941 404 -3349 410
rect -3283 444 -1691 450
rect -3283 410 -3271 444
rect -1703 410 -1691 444
rect -3283 404 -1691 410
rect -1625 444 -33 450
rect -1625 410 -1613 444
rect -45 410 -33 444
rect -1625 404 -33 410
rect 33 444 1625 450
rect 33 410 45 444
rect 1613 410 1625 444
rect 33 404 1625 410
rect 1691 444 3283 450
rect 1691 410 1703 444
rect 3271 410 3283 444
rect 1691 404 3283 410
rect 3349 444 4941 450
rect 3349 410 3361 444
rect 4929 410 4941 444
rect 3349 404 4941 410
rect -4997 314 -4951 326
rect -4997 254 -4991 314
rect -4957 254 -4951 314
rect -4997 242 -4951 254
rect -3339 314 -3293 326
rect -3339 254 -3333 314
rect -3299 254 -3293 314
rect -3339 242 -3293 254
rect -1681 314 -1635 326
rect -1681 254 -1675 314
rect -1641 254 -1635 314
rect -1681 242 -1635 254
rect -23 314 23 326
rect -23 254 -17 314
rect 17 254 23 314
rect -23 242 23 254
rect 1635 314 1681 326
rect 1635 254 1641 314
rect 1675 254 1681 314
rect 1635 242 1681 254
rect 3293 314 3339 326
rect 3293 254 3299 314
rect 3333 254 3339 314
rect 3293 242 3339 254
rect 4951 314 4997 326
rect 4951 254 4957 314
rect 4991 254 4997 314
rect 4951 242 4997 254
rect -4941 195 -3349 201
rect -4941 161 -4929 195
rect -3361 161 -3349 195
rect -4941 155 -3349 161
rect -3283 195 -1691 201
rect -3283 161 -3271 195
rect -1703 161 -1691 195
rect -3283 155 -1691 161
rect -1625 195 -33 201
rect -1625 161 -1613 195
rect -45 161 -33 195
rect -1625 155 -33 161
rect 33 195 1625 201
rect 33 161 45 195
rect 1613 161 1625 195
rect 33 155 1625 161
rect 1691 195 3283 201
rect 1691 161 1703 195
rect 3271 161 3283 195
rect 1691 155 3283 161
rect 3349 195 4941 201
rect 3349 161 3361 195
rect 4929 161 4941 195
rect 3349 155 4941 161
rect -4997 65 -4951 77
rect -4997 5 -4991 65
rect -4957 5 -4951 65
rect -4997 -7 -4951 5
rect -3339 65 -3293 77
rect -3339 5 -3333 65
rect -3299 5 -3293 65
rect -3339 -7 -3293 5
rect -1681 65 -1635 77
rect -1681 5 -1675 65
rect -1641 5 -1635 65
rect -1681 -7 -1635 5
rect -23 65 23 77
rect -23 5 -17 65
rect 17 5 23 65
rect -23 -7 23 5
rect 1635 65 1681 77
rect 1635 5 1641 65
rect 1675 5 1681 65
rect 1635 -7 1681 5
rect 3293 65 3339 77
rect 3293 5 3299 65
rect 3333 5 3339 65
rect 3293 -7 3339 5
rect 4951 65 4997 77
rect 4951 5 4957 65
rect 4991 5 4997 65
rect 4951 -7 4997 5
rect -4941 -54 -3349 -48
rect -4941 -88 -4929 -54
rect -3361 -88 -3349 -54
rect -4941 -94 -3349 -88
rect -3283 -54 -1691 -48
rect -3283 -88 -3271 -54
rect -1703 -88 -1691 -54
rect -3283 -94 -1691 -88
rect -1625 -54 -33 -48
rect -1625 -88 -1613 -54
rect -45 -88 -33 -54
rect -1625 -94 -33 -88
rect 33 -54 1625 -48
rect 33 -88 45 -54
rect 1613 -88 1625 -54
rect 33 -94 1625 -88
rect 1691 -54 3283 -48
rect 1691 -88 1703 -54
rect 3271 -88 3283 -54
rect 1691 -94 3283 -88
rect 3349 -54 4941 -48
rect 3349 -88 3361 -54
rect 4929 -88 4941 -54
rect 3349 -94 4941 -88
rect -4997 -184 -4951 -172
rect -4997 -244 -4991 -184
rect -4957 -244 -4951 -184
rect -4997 -256 -4951 -244
rect -3339 -184 -3293 -172
rect -3339 -244 -3333 -184
rect -3299 -244 -3293 -184
rect -3339 -256 -3293 -244
rect -1681 -184 -1635 -172
rect -1681 -244 -1675 -184
rect -1641 -244 -1635 -184
rect -1681 -256 -1635 -244
rect -23 -184 23 -172
rect -23 -244 -17 -184
rect 17 -244 23 -184
rect -23 -256 23 -244
rect 1635 -184 1681 -172
rect 1635 -244 1641 -184
rect 1675 -244 1681 -184
rect 1635 -256 1681 -244
rect 3293 -184 3339 -172
rect 3293 -244 3299 -184
rect 3333 -244 3339 -184
rect 3293 -256 3339 -244
rect 4951 -184 4997 -172
rect 4951 -244 4957 -184
rect 4991 -244 4997 -184
rect 4951 -256 4997 -244
rect -4941 -303 -3349 -297
rect -4941 -337 -4929 -303
rect -3361 -337 -3349 -303
rect -4941 -343 -3349 -337
rect -3283 -303 -1691 -297
rect -3283 -337 -3271 -303
rect -1703 -337 -1691 -303
rect -3283 -343 -1691 -337
rect -1625 -303 -33 -297
rect -1625 -337 -1613 -303
rect -45 -337 -33 -303
rect -1625 -343 -33 -337
rect 33 -303 1625 -297
rect 33 -337 45 -303
rect 1613 -337 1625 -303
rect 33 -343 1625 -337
rect 1691 -303 3283 -297
rect 1691 -337 1703 -303
rect 3271 -337 3283 -303
rect 1691 -343 3283 -337
rect 3349 -303 4941 -297
rect 3349 -337 3361 -303
rect 4929 -337 4941 -303
rect 3349 -343 4941 -337
rect -4997 -433 -4951 -421
rect -4997 -493 -4991 -433
rect -4957 -493 -4951 -433
rect -4997 -505 -4951 -493
rect -3339 -433 -3293 -421
rect -3339 -493 -3333 -433
rect -3299 -493 -3293 -433
rect -3339 -505 -3293 -493
rect -1681 -433 -1635 -421
rect -1681 -493 -1675 -433
rect -1641 -493 -1635 -433
rect -1681 -505 -1635 -493
rect -23 -433 23 -421
rect -23 -493 -17 -433
rect 17 -493 23 -433
rect -23 -505 23 -493
rect 1635 -433 1681 -421
rect 1635 -493 1641 -433
rect 1675 -493 1681 -433
rect 1635 -505 1681 -493
rect 3293 -433 3339 -421
rect 3293 -493 3299 -433
rect 3333 -493 3339 -433
rect 3293 -505 3339 -493
rect 4951 -433 4997 -421
rect 4951 -493 4957 -433
rect 4991 -493 4997 -433
rect 4951 -505 4997 -493
rect -4941 -552 -3349 -546
rect -4941 -586 -4929 -552
rect -3361 -586 -3349 -552
rect -4941 -592 -3349 -586
rect -3283 -552 -1691 -546
rect -3283 -586 -3271 -552
rect -1703 -586 -1691 -552
rect -3283 -592 -1691 -586
rect -1625 -552 -33 -546
rect -1625 -586 -1613 -552
rect -45 -586 -33 -552
rect -1625 -592 -33 -586
rect 33 -552 1625 -546
rect 33 -586 45 -552
rect 1613 -586 1625 -552
rect 33 -592 1625 -586
rect 1691 -552 3283 -546
rect 1691 -586 1703 -552
rect 3271 -586 3283 -552
rect 1691 -592 3283 -586
rect 3349 -552 4941 -546
rect 3349 -586 3361 -552
rect 4929 -586 4941 -552
rect 3349 -592 4941 -586
rect -4997 -682 -4951 -670
rect -4997 -742 -4991 -682
rect -4957 -742 -4951 -682
rect -4997 -754 -4951 -742
rect -3339 -682 -3293 -670
rect -3339 -742 -3333 -682
rect -3299 -742 -3293 -682
rect -3339 -754 -3293 -742
rect -1681 -682 -1635 -670
rect -1681 -742 -1675 -682
rect -1641 -742 -1635 -682
rect -1681 -754 -1635 -742
rect -23 -682 23 -670
rect -23 -742 -17 -682
rect 17 -742 23 -682
rect -23 -754 23 -742
rect 1635 -682 1681 -670
rect 1635 -742 1641 -682
rect 1675 -742 1681 -682
rect 1635 -754 1681 -742
rect 3293 -682 3339 -670
rect 3293 -742 3299 -682
rect 3333 -742 3339 -682
rect 3293 -754 3339 -742
rect 4951 -682 4997 -670
rect 4951 -742 4957 -682
rect 4991 -742 4997 -682
rect 4951 -754 4997 -742
rect -4941 -801 -3349 -795
rect -4941 -835 -4929 -801
rect -3361 -835 -3349 -801
rect -4941 -841 -3349 -835
rect -3283 -801 -1691 -795
rect -3283 -835 -3271 -801
rect -1703 -835 -1691 -801
rect -3283 -841 -1691 -835
rect -1625 -801 -33 -795
rect -1625 -835 -1613 -801
rect -45 -835 -33 -801
rect -1625 -841 -33 -835
rect 33 -801 1625 -795
rect 33 -835 45 -801
rect 1613 -835 1625 -801
rect 33 -841 1625 -835
rect 1691 -801 3283 -795
rect 1691 -835 1703 -801
rect 3271 -835 3283 -801
rect 1691 -841 3283 -835
rect 3349 -801 4941 -795
rect 3349 -835 3361 -801
rect 4929 -835 4941 -801
rect 3349 -841 4941 -835
rect -4997 -931 -4951 -919
rect -4997 -991 -4991 -931
rect -4957 -991 -4951 -931
rect -4997 -1003 -4951 -991
rect -3339 -931 -3293 -919
rect -3339 -991 -3333 -931
rect -3299 -991 -3293 -931
rect -3339 -1003 -3293 -991
rect -1681 -931 -1635 -919
rect -1681 -991 -1675 -931
rect -1641 -991 -1635 -931
rect -1681 -1003 -1635 -991
rect -23 -931 23 -919
rect -23 -991 -17 -931
rect 17 -991 23 -931
rect -23 -1003 23 -991
rect 1635 -931 1681 -919
rect 1635 -991 1641 -931
rect 1675 -991 1681 -931
rect 1635 -1003 1681 -991
rect 3293 -931 3339 -919
rect 3293 -991 3299 -931
rect 3333 -991 3339 -931
rect 3293 -1003 3339 -991
rect 4951 -931 4997 -919
rect 4951 -991 4957 -931
rect 4991 -991 4997 -931
rect 4951 -1003 4997 -991
rect -4941 -1050 -3349 -1044
rect -4941 -1084 -4929 -1050
rect -3361 -1084 -3349 -1050
rect -4941 -1090 -3349 -1084
rect -3283 -1050 -1691 -1044
rect -3283 -1084 -3271 -1050
rect -1703 -1084 -1691 -1050
rect -3283 -1090 -1691 -1084
rect -1625 -1050 -33 -1044
rect -1625 -1084 -1613 -1050
rect -45 -1084 -33 -1050
rect -1625 -1090 -33 -1084
rect 33 -1050 1625 -1044
rect 33 -1084 45 -1050
rect 1613 -1084 1625 -1050
rect 33 -1090 1625 -1084
rect 1691 -1050 3283 -1044
rect 1691 -1084 1703 -1050
rect 3271 -1084 3283 -1050
rect 1691 -1090 3283 -1084
rect 3349 -1050 4941 -1044
rect 3349 -1084 3361 -1050
rect 4929 -1084 4941 -1050
rect 3349 -1090 4941 -1084
<< properties >>
string FIXED_BBOX -5108 -1205 5108 1205
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 8 m 9 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
