magic
tech sky130A
magscale 1 2
timestamp 1712153244
<< nwell >>
rect -20026 -2405 20026 2405
<< mvnsubdiff >>
rect -19960 2327 19960 2339
rect -19960 2293 -19852 2327
rect 19852 2293 19960 2327
rect -19960 2281 19960 2293
rect -19960 2231 -19902 2281
rect -19960 -2231 -19948 2231
rect -19914 -2231 -19902 2231
rect 19902 2231 19960 2281
rect -19960 -2281 -19902 -2231
rect 19902 -2231 19914 2231
rect 19948 -2231 19960 2231
rect 19902 -2281 19960 -2231
rect -19960 -2293 19960 -2281
rect -19960 -2327 -19852 -2293
rect 19852 -2327 19960 -2293
rect -19960 -2339 19960 -2327
<< mvnsubdiffcont >>
rect -19852 2293 19852 2327
rect -19948 -2231 -19914 2231
rect 19914 -2231 19948 2231
rect -19852 -2327 19852 -2293
<< xpolycontact >>
rect -19797 1744 -19515 2176
rect -19797 -2176 -19515 -1744
rect -19419 1744 -19137 2176
rect -19419 -2176 -19137 -1744
rect -19041 1744 -18759 2176
rect -19041 -2176 -18759 -1744
rect -18663 1744 -18381 2176
rect -18663 -2176 -18381 -1744
rect -18285 1744 -18003 2176
rect -18285 -2176 -18003 -1744
rect -17907 1744 -17625 2176
rect -17907 -2176 -17625 -1744
rect -17529 1744 -17247 2176
rect -17529 -2176 -17247 -1744
rect -17151 1744 -16869 2176
rect -17151 -2176 -16869 -1744
rect -16773 1744 -16491 2176
rect -16773 -2176 -16491 -1744
rect -16395 1744 -16113 2176
rect -16395 -2176 -16113 -1744
rect -16017 1744 -15735 2176
rect -16017 -2176 -15735 -1744
rect -15639 1744 -15357 2176
rect -15639 -2176 -15357 -1744
rect -15261 1744 -14979 2176
rect -15261 -2176 -14979 -1744
rect -14883 1744 -14601 2176
rect -14883 -2176 -14601 -1744
rect -14505 1744 -14223 2176
rect -14505 -2176 -14223 -1744
rect -14127 1744 -13845 2176
rect -14127 -2176 -13845 -1744
rect -13749 1744 -13467 2176
rect -13749 -2176 -13467 -1744
rect -13371 1744 -13089 2176
rect -13371 -2176 -13089 -1744
rect -12993 1744 -12711 2176
rect -12993 -2176 -12711 -1744
rect -12615 1744 -12333 2176
rect -12615 -2176 -12333 -1744
rect -12237 1744 -11955 2176
rect -12237 -2176 -11955 -1744
rect -11859 1744 -11577 2176
rect -11859 -2176 -11577 -1744
rect -11481 1744 -11199 2176
rect -11481 -2176 -11199 -1744
rect -11103 1744 -10821 2176
rect -11103 -2176 -10821 -1744
rect -10725 1744 -10443 2176
rect -10725 -2176 -10443 -1744
rect -10347 1744 -10065 2176
rect -10347 -2176 -10065 -1744
rect -9969 1744 -9687 2176
rect -9969 -2176 -9687 -1744
rect -9591 1744 -9309 2176
rect -9591 -2176 -9309 -1744
rect -9213 1744 -8931 2176
rect -9213 -2176 -8931 -1744
rect -8835 1744 -8553 2176
rect -8835 -2176 -8553 -1744
rect -8457 1744 -8175 2176
rect -8457 -2176 -8175 -1744
rect -8079 1744 -7797 2176
rect -8079 -2176 -7797 -1744
rect -7701 1744 -7419 2176
rect -7701 -2176 -7419 -1744
rect -7323 1744 -7041 2176
rect -7323 -2176 -7041 -1744
rect -6945 1744 -6663 2176
rect -6945 -2176 -6663 -1744
rect -6567 1744 -6285 2176
rect -6567 -2176 -6285 -1744
rect -6189 1744 -5907 2176
rect -6189 -2176 -5907 -1744
rect -5811 1744 -5529 2176
rect -5811 -2176 -5529 -1744
rect -5433 1744 -5151 2176
rect -5433 -2176 -5151 -1744
rect -5055 1744 -4773 2176
rect -5055 -2176 -4773 -1744
rect -4677 1744 -4395 2176
rect -4677 -2176 -4395 -1744
rect -4299 1744 -4017 2176
rect -4299 -2176 -4017 -1744
rect -3921 1744 -3639 2176
rect -3921 -2176 -3639 -1744
rect -3543 1744 -3261 2176
rect -3543 -2176 -3261 -1744
rect -3165 1744 -2883 2176
rect -3165 -2176 -2883 -1744
rect -2787 1744 -2505 2176
rect -2787 -2176 -2505 -1744
rect -2409 1744 -2127 2176
rect -2409 -2176 -2127 -1744
rect -2031 1744 -1749 2176
rect -2031 -2176 -1749 -1744
rect -1653 1744 -1371 2176
rect -1653 -2176 -1371 -1744
rect -1275 1744 -993 2176
rect -1275 -2176 -993 -1744
rect -897 1744 -615 2176
rect -897 -2176 -615 -1744
rect -519 1744 -237 2176
rect -519 -2176 -237 -1744
rect -141 1744 141 2176
rect -141 -2176 141 -1744
rect 237 1744 519 2176
rect 237 -2176 519 -1744
rect 615 1744 897 2176
rect 615 -2176 897 -1744
rect 993 1744 1275 2176
rect 993 -2176 1275 -1744
rect 1371 1744 1653 2176
rect 1371 -2176 1653 -1744
rect 1749 1744 2031 2176
rect 1749 -2176 2031 -1744
rect 2127 1744 2409 2176
rect 2127 -2176 2409 -1744
rect 2505 1744 2787 2176
rect 2505 -2176 2787 -1744
rect 2883 1744 3165 2176
rect 2883 -2176 3165 -1744
rect 3261 1744 3543 2176
rect 3261 -2176 3543 -1744
rect 3639 1744 3921 2176
rect 3639 -2176 3921 -1744
rect 4017 1744 4299 2176
rect 4017 -2176 4299 -1744
rect 4395 1744 4677 2176
rect 4395 -2176 4677 -1744
rect 4773 1744 5055 2176
rect 4773 -2176 5055 -1744
rect 5151 1744 5433 2176
rect 5151 -2176 5433 -1744
rect 5529 1744 5811 2176
rect 5529 -2176 5811 -1744
rect 5907 1744 6189 2176
rect 5907 -2176 6189 -1744
rect 6285 1744 6567 2176
rect 6285 -2176 6567 -1744
rect 6663 1744 6945 2176
rect 6663 -2176 6945 -1744
rect 7041 1744 7323 2176
rect 7041 -2176 7323 -1744
rect 7419 1744 7701 2176
rect 7419 -2176 7701 -1744
rect 7797 1744 8079 2176
rect 7797 -2176 8079 -1744
rect 8175 1744 8457 2176
rect 8175 -2176 8457 -1744
rect 8553 1744 8835 2176
rect 8553 -2176 8835 -1744
rect 8931 1744 9213 2176
rect 8931 -2176 9213 -1744
rect 9309 1744 9591 2176
rect 9309 -2176 9591 -1744
rect 9687 1744 9969 2176
rect 9687 -2176 9969 -1744
rect 10065 1744 10347 2176
rect 10065 -2176 10347 -1744
rect 10443 1744 10725 2176
rect 10443 -2176 10725 -1744
rect 10821 1744 11103 2176
rect 10821 -2176 11103 -1744
rect 11199 1744 11481 2176
rect 11199 -2176 11481 -1744
rect 11577 1744 11859 2176
rect 11577 -2176 11859 -1744
rect 11955 1744 12237 2176
rect 11955 -2176 12237 -1744
rect 12333 1744 12615 2176
rect 12333 -2176 12615 -1744
rect 12711 1744 12993 2176
rect 12711 -2176 12993 -1744
rect 13089 1744 13371 2176
rect 13089 -2176 13371 -1744
rect 13467 1744 13749 2176
rect 13467 -2176 13749 -1744
rect 13845 1744 14127 2176
rect 13845 -2176 14127 -1744
rect 14223 1744 14505 2176
rect 14223 -2176 14505 -1744
rect 14601 1744 14883 2176
rect 14601 -2176 14883 -1744
rect 14979 1744 15261 2176
rect 14979 -2176 15261 -1744
rect 15357 1744 15639 2176
rect 15357 -2176 15639 -1744
rect 15735 1744 16017 2176
rect 15735 -2176 16017 -1744
rect 16113 1744 16395 2176
rect 16113 -2176 16395 -1744
rect 16491 1744 16773 2176
rect 16491 -2176 16773 -1744
rect 16869 1744 17151 2176
rect 16869 -2176 17151 -1744
rect 17247 1744 17529 2176
rect 17247 -2176 17529 -1744
rect 17625 1744 17907 2176
rect 17625 -2176 17907 -1744
rect 18003 1744 18285 2176
rect 18003 -2176 18285 -1744
rect 18381 1744 18663 2176
rect 18381 -2176 18663 -1744
rect 18759 1744 19041 2176
rect 18759 -2176 19041 -1744
rect 19137 1744 19419 2176
rect 19137 -2176 19419 -1744
rect 19515 1744 19797 2176
rect 19515 -2176 19797 -1744
<< xpolyres >>
rect -19797 -1744 -19515 1744
rect -19419 -1744 -19137 1744
rect -19041 -1744 -18759 1744
rect -18663 -1744 -18381 1744
rect -18285 -1744 -18003 1744
rect -17907 -1744 -17625 1744
rect -17529 -1744 -17247 1744
rect -17151 -1744 -16869 1744
rect -16773 -1744 -16491 1744
rect -16395 -1744 -16113 1744
rect -16017 -1744 -15735 1744
rect -15639 -1744 -15357 1744
rect -15261 -1744 -14979 1744
rect -14883 -1744 -14601 1744
rect -14505 -1744 -14223 1744
rect -14127 -1744 -13845 1744
rect -13749 -1744 -13467 1744
rect -13371 -1744 -13089 1744
rect -12993 -1744 -12711 1744
rect -12615 -1744 -12333 1744
rect -12237 -1744 -11955 1744
rect -11859 -1744 -11577 1744
rect -11481 -1744 -11199 1744
rect -11103 -1744 -10821 1744
rect -10725 -1744 -10443 1744
rect -10347 -1744 -10065 1744
rect -9969 -1744 -9687 1744
rect -9591 -1744 -9309 1744
rect -9213 -1744 -8931 1744
rect -8835 -1744 -8553 1744
rect -8457 -1744 -8175 1744
rect -8079 -1744 -7797 1744
rect -7701 -1744 -7419 1744
rect -7323 -1744 -7041 1744
rect -6945 -1744 -6663 1744
rect -6567 -1744 -6285 1744
rect -6189 -1744 -5907 1744
rect -5811 -1744 -5529 1744
rect -5433 -1744 -5151 1744
rect -5055 -1744 -4773 1744
rect -4677 -1744 -4395 1744
rect -4299 -1744 -4017 1744
rect -3921 -1744 -3639 1744
rect -3543 -1744 -3261 1744
rect -3165 -1744 -2883 1744
rect -2787 -1744 -2505 1744
rect -2409 -1744 -2127 1744
rect -2031 -1744 -1749 1744
rect -1653 -1744 -1371 1744
rect -1275 -1744 -993 1744
rect -897 -1744 -615 1744
rect -519 -1744 -237 1744
rect -141 -1744 141 1744
rect 237 -1744 519 1744
rect 615 -1744 897 1744
rect 993 -1744 1275 1744
rect 1371 -1744 1653 1744
rect 1749 -1744 2031 1744
rect 2127 -1744 2409 1744
rect 2505 -1744 2787 1744
rect 2883 -1744 3165 1744
rect 3261 -1744 3543 1744
rect 3639 -1744 3921 1744
rect 4017 -1744 4299 1744
rect 4395 -1744 4677 1744
rect 4773 -1744 5055 1744
rect 5151 -1744 5433 1744
rect 5529 -1744 5811 1744
rect 5907 -1744 6189 1744
rect 6285 -1744 6567 1744
rect 6663 -1744 6945 1744
rect 7041 -1744 7323 1744
rect 7419 -1744 7701 1744
rect 7797 -1744 8079 1744
rect 8175 -1744 8457 1744
rect 8553 -1744 8835 1744
rect 8931 -1744 9213 1744
rect 9309 -1744 9591 1744
rect 9687 -1744 9969 1744
rect 10065 -1744 10347 1744
rect 10443 -1744 10725 1744
rect 10821 -1744 11103 1744
rect 11199 -1744 11481 1744
rect 11577 -1744 11859 1744
rect 11955 -1744 12237 1744
rect 12333 -1744 12615 1744
rect 12711 -1744 12993 1744
rect 13089 -1744 13371 1744
rect 13467 -1744 13749 1744
rect 13845 -1744 14127 1744
rect 14223 -1744 14505 1744
rect 14601 -1744 14883 1744
rect 14979 -1744 15261 1744
rect 15357 -1744 15639 1744
rect 15735 -1744 16017 1744
rect 16113 -1744 16395 1744
rect 16491 -1744 16773 1744
rect 16869 -1744 17151 1744
rect 17247 -1744 17529 1744
rect 17625 -1744 17907 1744
rect 18003 -1744 18285 1744
rect 18381 -1744 18663 1744
rect 18759 -1744 19041 1744
rect 19137 -1744 19419 1744
rect 19515 -1744 19797 1744
<< locali >>
rect -19948 2293 -19852 2327
rect 19852 2293 19948 2327
rect -19948 2231 -19914 2293
rect 19914 2231 19948 2293
rect -19948 -2293 -19914 -2231
rect 19914 -2293 19948 -2231
rect -19948 -2327 -19852 -2293
rect 19852 -2327 19948 -2293
<< viali >>
rect -19781 1761 -19531 2158
rect -19403 1761 -19153 2158
rect -19025 1761 -18775 2158
rect -18647 1761 -18397 2158
rect -18269 1761 -18019 2158
rect -17891 1761 -17641 2158
rect -17513 1761 -17263 2158
rect -17135 1761 -16885 2158
rect -16757 1761 -16507 2158
rect -16379 1761 -16129 2158
rect -16001 1761 -15751 2158
rect -15623 1761 -15373 2158
rect -15245 1761 -14995 2158
rect -14867 1761 -14617 2158
rect -14489 1761 -14239 2158
rect -14111 1761 -13861 2158
rect -13733 1761 -13483 2158
rect -13355 1761 -13105 2158
rect -12977 1761 -12727 2158
rect -12599 1761 -12349 2158
rect -12221 1761 -11971 2158
rect -11843 1761 -11593 2158
rect -11465 1761 -11215 2158
rect -11087 1761 -10837 2158
rect -10709 1761 -10459 2158
rect -10331 1761 -10081 2158
rect -9953 1761 -9703 2158
rect -9575 1761 -9325 2158
rect -9197 1761 -8947 2158
rect -8819 1761 -8569 2158
rect -8441 1761 -8191 2158
rect -8063 1761 -7813 2158
rect -7685 1761 -7435 2158
rect -7307 1761 -7057 2158
rect -6929 1761 -6679 2158
rect -6551 1761 -6301 2158
rect -6173 1761 -5923 2158
rect -5795 1761 -5545 2158
rect -5417 1761 -5167 2158
rect -5039 1761 -4789 2158
rect -4661 1761 -4411 2158
rect -4283 1761 -4033 2158
rect -3905 1761 -3655 2158
rect -3527 1761 -3277 2158
rect -3149 1761 -2899 2158
rect -2771 1761 -2521 2158
rect -2393 1761 -2143 2158
rect -2015 1761 -1765 2158
rect -1637 1761 -1387 2158
rect -1259 1761 -1009 2158
rect -881 1761 -631 2158
rect -503 1761 -253 2158
rect -125 1761 125 2158
rect 253 1761 503 2158
rect 631 1761 881 2158
rect 1009 1761 1259 2158
rect 1387 1761 1637 2158
rect 1765 1761 2015 2158
rect 2143 1761 2393 2158
rect 2521 1761 2771 2158
rect 2899 1761 3149 2158
rect 3277 1761 3527 2158
rect 3655 1761 3905 2158
rect 4033 1761 4283 2158
rect 4411 1761 4661 2158
rect 4789 1761 5039 2158
rect 5167 1761 5417 2158
rect 5545 1761 5795 2158
rect 5923 1761 6173 2158
rect 6301 1761 6551 2158
rect 6679 1761 6929 2158
rect 7057 1761 7307 2158
rect 7435 1761 7685 2158
rect 7813 1761 8063 2158
rect 8191 1761 8441 2158
rect 8569 1761 8819 2158
rect 8947 1761 9197 2158
rect 9325 1761 9575 2158
rect 9703 1761 9953 2158
rect 10081 1761 10331 2158
rect 10459 1761 10709 2158
rect 10837 1761 11087 2158
rect 11215 1761 11465 2158
rect 11593 1761 11843 2158
rect 11971 1761 12221 2158
rect 12349 1761 12599 2158
rect 12727 1761 12977 2158
rect 13105 1761 13355 2158
rect 13483 1761 13733 2158
rect 13861 1761 14111 2158
rect 14239 1761 14489 2158
rect 14617 1761 14867 2158
rect 14995 1761 15245 2158
rect 15373 1761 15623 2158
rect 15751 1761 16001 2158
rect 16129 1761 16379 2158
rect 16507 1761 16757 2158
rect 16885 1761 17135 2158
rect 17263 1761 17513 2158
rect 17641 1761 17891 2158
rect 18019 1761 18269 2158
rect 18397 1761 18647 2158
rect 18775 1761 19025 2158
rect 19153 1761 19403 2158
rect 19531 1761 19781 2158
rect -19781 -2158 -19531 -1761
rect -19403 -2158 -19153 -1761
rect -19025 -2158 -18775 -1761
rect -18647 -2158 -18397 -1761
rect -18269 -2158 -18019 -1761
rect -17891 -2158 -17641 -1761
rect -17513 -2158 -17263 -1761
rect -17135 -2158 -16885 -1761
rect -16757 -2158 -16507 -1761
rect -16379 -2158 -16129 -1761
rect -16001 -2158 -15751 -1761
rect -15623 -2158 -15373 -1761
rect -15245 -2158 -14995 -1761
rect -14867 -2158 -14617 -1761
rect -14489 -2158 -14239 -1761
rect -14111 -2158 -13861 -1761
rect -13733 -2158 -13483 -1761
rect -13355 -2158 -13105 -1761
rect -12977 -2158 -12727 -1761
rect -12599 -2158 -12349 -1761
rect -12221 -2158 -11971 -1761
rect -11843 -2158 -11593 -1761
rect -11465 -2158 -11215 -1761
rect -11087 -2158 -10837 -1761
rect -10709 -2158 -10459 -1761
rect -10331 -2158 -10081 -1761
rect -9953 -2158 -9703 -1761
rect -9575 -2158 -9325 -1761
rect -9197 -2158 -8947 -1761
rect -8819 -2158 -8569 -1761
rect -8441 -2158 -8191 -1761
rect -8063 -2158 -7813 -1761
rect -7685 -2158 -7435 -1761
rect -7307 -2158 -7057 -1761
rect -6929 -2158 -6679 -1761
rect -6551 -2158 -6301 -1761
rect -6173 -2158 -5923 -1761
rect -5795 -2158 -5545 -1761
rect -5417 -2158 -5167 -1761
rect -5039 -2158 -4789 -1761
rect -4661 -2158 -4411 -1761
rect -4283 -2158 -4033 -1761
rect -3905 -2158 -3655 -1761
rect -3527 -2158 -3277 -1761
rect -3149 -2158 -2899 -1761
rect -2771 -2158 -2521 -1761
rect -2393 -2158 -2143 -1761
rect -2015 -2158 -1765 -1761
rect -1637 -2158 -1387 -1761
rect -1259 -2158 -1009 -1761
rect -881 -2158 -631 -1761
rect -503 -2158 -253 -1761
rect -125 -2158 125 -1761
rect 253 -2158 503 -1761
rect 631 -2158 881 -1761
rect 1009 -2158 1259 -1761
rect 1387 -2158 1637 -1761
rect 1765 -2158 2015 -1761
rect 2143 -2158 2393 -1761
rect 2521 -2158 2771 -1761
rect 2899 -2158 3149 -1761
rect 3277 -2158 3527 -1761
rect 3655 -2158 3905 -1761
rect 4033 -2158 4283 -1761
rect 4411 -2158 4661 -1761
rect 4789 -2158 5039 -1761
rect 5167 -2158 5417 -1761
rect 5545 -2158 5795 -1761
rect 5923 -2158 6173 -1761
rect 6301 -2158 6551 -1761
rect 6679 -2158 6929 -1761
rect 7057 -2158 7307 -1761
rect 7435 -2158 7685 -1761
rect 7813 -2158 8063 -1761
rect 8191 -2158 8441 -1761
rect 8569 -2158 8819 -1761
rect 8947 -2158 9197 -1761
rect 9325 -2158 9575 -1761
rect 9703 -2158 9953 -1761
rect 10081 -2158 10331 -1761
rect 10459 -2158 10709 -1761
rect 10837 -2158 11087 -1761
rect 11215 -2158 11465 -1761
rect 11593 -2158 11843 -1761
rect 11971 -2158 12221 -1761
rect 12349 -2158 12599 -1761
rect 12727 -2158 12977 -1761
rect 13105 -2158 13355 -1761
rect 13483 -2158 13733 -1761
rect 13861 -2158 14111 -1761
rect 14239 -2158 14489 -1761
rect 14617 -2158 14867 -1761
rect 14995 -2158 15245 -1761
rect 15373 -2158 15623 -1761
rect 15751 -2158 16001 -1761
rect 16129 -2158 16379 -1761
rect 16507 -2158 16757 -1761
rect 16885 -2158 17135 -1761
rect 17263 -2158 17513 -1761
rect 17641 -2158 17891 -1761
rect 18019 -2158 18269 -1761
rect 18397 -2158 18647 -1761
rect 18775 -2158 19025 -1761
rect 19153 -2158 19403 -1761
rect 19531 -2158 19781 -1761
<< metal1 >>
rect -19787 2158 -19525 2170
rect -19787 1761 -19781 2158
rect -19531 1761 -19525 2158
rect -19787 1749 -19525 1761
rect -19409 2158 -19147 2170
rect -19409 1761 -19403 2158
rect -19153 1761 -19147 2158
rect -19409 1749 -19147 1761
rect -19031 2158 -18769 2170
rect -19031 1761 -19025 2158
rect -18775 1761 -18769 2158
rect -19031 1749 -18769 1761
rect -18653 2158 -18391 2170
rect -18653 1761 -18647 2158
rect -18397 1761 -18391 2158
rect -18653 1749 -18391 1761
rect -18275 2158 -18013 2170
rect -18275 1761 -18269 2158
rect -18019 1761 -18013 2158
rect -18275 1749 -18013 1761
rect -17897 2158 -17635 2170
rect -17897 1761 -17891 2158
rect -17641 1761 -17635 2158
rect -17897 1749 -17635 1761
rect -17519 2158 -17257 2170
rect -17519 1761 -17513 2158
rect -17263 1761 -17257 2158
rect -17519 1749 -17257 1761
rect -17141 2158 -16879 2170
rect -17141 1761 -17135 2158
rect -16885 1761 -16879 2158
rect -17141 1749 -16879 1761
rect -16763 2158 -16501 2170
rect -16763 1761 -16757 2158
rect -16507 1761 -16501 2158
rect -16763 1749 -16501 1761
rect -16385 2158 -16123 2170
rect -16385 1761 -16379 2158
rect -16129 1761 -16123 2158
rect -16385 1749 -16123 1761
rect -16007 2158 -15745 2170
rect -16007 1761 -16001 2158
rect -15751 1761 -15745 2158
rect -16007 1749 -15745 1761
rect -15629 2158 -15367 2170
rect -15629 1761 -15623 2158
rect -15373 1761 -15367 2158
rect -15629 1749 -15367 1761
rect -15251 2158 -14989 2170
rect -15251 1761 -15245 2158
rect -14995 1761 -14989 2158
rect -15251 1749 -14989 1761
rect -14873 2158 -14611 2170
rect -14873 1761 -14867 2158
rect -14617 1761 -14611 2158
rect -14873 1749 -14611 1761
rect -14495 2158 -14233 2170
rect -14495 1761 -14489 2158
rect -14239 1761 -14233 2158
rect -14495 1749 -14233 1761
rect -14117 2158 -13855 2170
rect -14117 1761 -14111 2158
rect -13861 1761 -13855 2158
rect -14117 1749 -13855 1761
rect -13739 2158 -13477 2170
rect -13739 1761 -13733 2158
rect -13483 1761 -13477 2158
rect -13739 1749 -13477 1761
rect -13361 2158 -13099 2170
rect -13361 1761 -13355 2158
rect -13105 1761 -13099 2158
rect -13361 1749 -13099 1761
rect -12983 2158 -12721 2170
rect -12983 1761 -12977 2158
rect -12727 1761 -12721 2158
rect -12983 1749 -12721 1761
rect -12605 2158 -12343 2170
rect -12605 1761 -12599 2158
rect -12349 1761 -12343 2158
rect -12605 1749 -12343 1761
rect -12227 2158 -11965 2170
rect -12227 1761 -12221 2158
rect -11971 1761 -11965 2158
rect -12227 1749 -11965 1761
rect -11849 2158 -11587 2170
rect -11849 1761 -11843 2158
rect -11593 1761 -11587 2158
rect -11849 1749 -11587 1761
rect -11471 2158 -11209 2170
rect -11471 1761 -11465 2158
rect -11215 1761 -11209 2158
rect -11471 1749 -11209 1761
rect -11093 2158 -10831 2170
rect -11093 1761 -11087 2158
rect -10837 1761 -10831 2158
rect -11093 1749 -10831 1761
rect -10715 2158 -10453 2170
rect -10715 1761 -10709 2158
rect -10459 1761 -10453 2158
rect -10715 1749 -10453 1761
rect -10337 2158 -10075 2170
rect -10337 1761 -10331 2158
rect -10081 1761 -10075 2158
rect -10337 1749 -10075 1761
rect -9959 2158 -9697 2170
rect -9959 1761 -9953 2158
rect -9703 1761 -9697 2158
rect -9959 1749 -9697 1761
rect -9581 2158 -9319 2170
rect -9581 1761 -9575 2158
rect -9325 1761 -9319 2158
rect -9581 1749 -9319 1761
rect -9203 2158 -8941 2170
rect -9203 1761 -9197 2158
rect -8947 1761 -8941 2158
rect -9203 1749 -8941 1761
rect -8825 2158 -8563 2170
rect -8825 1761 -8819 2158
rect -8569 1761 -8563 2158
rect -8825 1749 -8563 1761
rect -8447 2158 -8185 2170
rect -8447 1761 -8441 2158
rect -8191 1761 -8185 2158
rect -8447 1749 -8185 1761
rect -8069 2158 -7807 2170
rect -8069 1761 -8063 2158
rect -7813 1761 -7807 2158
rect -8069 1749 -7807 1761
rect -7691 2158 -7429 2170
rect -7691 1761 -7685 2158
rect -7435 1761 -7429 2158
rect -7691 1749 -7429 1761
rect -7313 2158 -7051 2170
rect -7313 1761 -7307 2158
rect -7057 1761 -7051 2158
rect -7313 1749 -7051 1761
rect -6935 2158 -6673 2170
rect -6935 1761 -6929 2158
rect -6679 1761 -6673 2158
rect -6935 1749 -6673 1761
rect -6557 2158 -6295 2170
rect -6557 1761 -6551 2158
rect -6301 1761 -6295 2158
rect -6557 1749 -6295 1761
rect -6179 2158 -5917 2170
rect -6179 1761 -6173 2158
rect -5923 1761 -5917 2158
rect -6179 1749 -5917 1761
rect -5801 2158 -5539 2170
rect -5801 1761 -5795 2158
rect -5545 1761 -5539 2158
rect -5801 1749 -5539 1761
rect -5423 2158 -5161 2170
rect -5423 1761 -5417 2158
rect -5167 1761 -5161 2158
rect -5423 1749 -5161 1761
rect -5045 2158 -4783 2170
rect -5045 1761 -5039 2158
rect -4789 1761 -4783 2158
rect -5045 1749 -4783 1761
rect -4667 2158 -4405 2170
rect -4667 1761 -4661 2158
rect -4411 1761 -4405 2158
rect -4667 1749 -4405 1761
rect -4289 2158 -4027 2170
rect -4289 1761 -4283 2158
rect -4033 1761 -4027 2158
rect -4289 1749 -4027 1761
rect -3911 2158 -3649 2170
rect -3911 1761 -3905 2158
rect -3655 1761 -3649 2158
rect -3911 1749 -3649 1761
rect -3533 2158 -3271 2170
rect -3533 1761 -3527 2158
rect -3277 1761 -3271 2158
rect -3533 1749 -3271 1761
rect -3155 2158 -2893 2170
rect -3155 1761 -3149 2158
rect -2899 1761 -2893 2158
rect -3155 1749 -2893 1761
rect -2777 2158 -2515 2170
rect -2777 1761 -2771 2158
rect -2521 1761 -2515 2158
rect -2777 1749 -2515 1761
rect -2399 2158 -2137 2170
rect -2399 1761 -2393 2158
rect -2143 1761 -2137 2158
rect -2399 1749 -2137 1761
rect -2021 2158 -1759 2170
rect -2021 1761 -2015 2158
rect -1765 1761 -1759 2158
rect -2021 1749 -1759 1761
rect -1643 2158 -1381 2170
rect -1643 1761 -1637 2158
rect -1387 1761 -1381 2158
rect -1643 1749 -1381 1761
rect -1265 2158 -1003 2170
rect -1265 1761 -1259 2158
rect -1009 1761 -1003 2158
rect -1265 1749 -1003 1761
rect -887 2158 -625 2170
rect -887 1761 -881 2158
rect -631 1761 -625 2158
rect -887 1749 -625 1761
rect -509 2158 -247 2170
rect -509 1761 -503 2158
rect -253 1761 -247 2158
rect -509 1749 -247 1761
rect -131 2158 131 2170
rect -131 1761 -125 2158
rect 125 1761 131 2158
rect -131 1749 131 1761
rect 247 2158 509 2170
rect 247 1761 253 2158
rect 503 1761 509 2158
rect 247 1749 509 1761
rect 625 2158 887 2170
rect 625 1761 631 2158
rect 881 1761 887 2158
rect 625 1749 887 1761
rect 1003 2158 1265 2170
rect 1003 1761 1009 2158
rect 1259 1761 1265 2158
rect 1003 1749 1265 1761
rect 1381 2158 1643 2170
rect 1381 1761 1387 2158
rect 1637 1761 1643 2158
rect 1381 1749 1643 1761
rect 1759 2158 2021 2170
rect 1759 1761 1765 2158
rect 2015 1761 2021 2158
rect 1759 1749 2021 1761
rect 2137 2158 2399 2170
rect 2137 1761 2143 2158
rect 2393 1761 2399 2158
rect 2137 1749 2399 1761
rect 2515 2158 2777 2170
rect 2515 1761 2521 2158
rect 2771 1761 2777 2158
rect 2515 1749 2777 1761
rect 2893 2158 3155 2170
rect 2893 1761 2899 2158
rect 3149 1761 3155 2158
rect 2893 1749 3155 1761
rect 3271 2158 3533 2170
rect 3271 1761 3277 2158
rect 3527 1761 3533 2158
rect 3271 1749 3533 1761
rect 3649 2158 3911 2170
rect 3649 1761 3655 2158
rect 3905 1761 3911 2158
rect 3649 1749 3911 1761
rect 4027 2158 4289 2170
rect 4027 1761 4033 2158
rect 4283 1761 4289 2158
rect 4027 1749 4289 1761
rect 4405 2158 4667 2170
rect 4405 1761 4411 2158
rect 4661 1761 4667 2158
rect 4405 1749 4667 1761
rect 4783 2158 5045 2170
rect 4783 1761 4789 2158
rect 5039 1761 5045 2158
rect 4783 1749 5045 1761
rect 5161 2158 5423 2170
rect 5161 1761 5167 2158
rect 5417 1761 5423 2158
rect 5161 1749 5423 1761
rect 5539 2158 5801 2170
rect 5539 1761 5545 2158
rect 5795 1761 5801 2158
rect 5539 1749 5801 1761
rect 5917 2158 6179 2170
rect 5917 1761 5923 2158
rect 6173 1761 6179 2158
rect 5917 1749 6179 1761
rect 6295 2158 6557 2170
rect 6295 1761 6301 2158
rect 6551 1761 6557 2158
rect 6295 1749 6557 1761
rect 6673 2158 6935 2170
rect 6673 1761 6679 2158
rect 6929 1761 6935 2158
rect 6673 1749 6935 1761
rect 7051 2158 7313 2170
rect 7051 1761 7057 2158
rect 7307 1761 7313 2158
rect 7051 1749 7313 1761
rect 7429 2158 7691 2170
rect 7429 1761 7435 2158
rect 7685 1761 7691 2158
rect 7429 1749 7691 1761
rect 7807 2158 8069 2170
rect 7807 1761 7813 2158
rect 8063 1761 8069 2158
rect 7807 1749 8069 1761
rect 8185 2158 8447 2170
rect 8185 1761 8191 2158
rect 8441 1761 8447 2158
rect 8185 1749 8447 1761
rect 8563 2158 8825 2170
rect 8563 1761 8569 2158
rect 8819 1761 8825 2158
rect 8563 1749 8825 1761
rect 8941 2158 9203 2170
rect 8941 1761 8947 2158
rect 9197 1761 9203 2158
rect 8941 1749 9203 1761
rect 9319 2158 9581 2170
rect 9319 1761 9325 2158
rect 9575 1761 9581 2158
rect 9319 1749 9581 1761
rect 9697 2158 9959 2170
rect 9697 1761 9703 2158
rect 9953 1761 9959 2158
rect 9697 1749 9959 1761
rect 10075 2158 10337 2170
rect 10075 1761 10081 2158
rect 10331 1761 10337 2158
rect 10075 1749 10337 1761
rect 10453 2158 10715 2170
rect 10453 1761 10459 2158
rect 10709 1761 10715 2158
rect 10453 1749 10715 1761
rect 10831 2158 11093 2170
rect 10831 1761 10837 2158
rect 11087 1761 11093 2158
rect 10831 1749 11093 1761
rect 11209 2158 11471 2170
rect 11209 1761 11215 2158
rect 11465 1761 11471 2158
rect 11209 1749 11471 1761
rect 11587 2158 11849 2170
rect 11587 1761 11593 2158
rect 11843 1761 11849 2158
rect 11587 1749 11849 1761
rect 11965 2158 12227 2170
rect 11965 1761 11971 2158
rect 12221 1761 12227 2158
rect 11965 1749 12227 1761
rect 12343 2158 12605 2170
rect 12343 1761 12349 2158
rect 12599 1761 12605 2158
rect 12343 1749 12605 1761
rect 12721 2158 12983 2170
rect 12721 1761 12727 2158
rect 12977 1761 12983 2158
rect 12721 1749 12983 1761
rect 13099 2158 13361 2170
rect 13099 1761 13105 2158
rect 13355 1761 13361 2158
rect 13099 1749 13361 1761
rect 13477 2158 13739 2170
rect 13477 1761 13483 2158
rect 13733 1761 13739 2158
rect 13477 1749 13739 1761
rect 13855 2158 14117 2170
rect 13855 1761 13861 2158
rect 14111 1761 14117 2158
rect 13855 1749 14117 1761
rect 14233 2158 14495 2170
rect 14233 1761 14239 2158
rect 14489 1761 14495 2158
rect 14233 1749 14495 1761
rect 14611 2158 14873 2170
rect 14611 1761 14617 2158
rect 14867 1761 14873 2158
rect 14611 1749 14873 1761
rect 14989 2158 15251 2170
rect 14989 1761 14995 2158
rect 15245 1761 15251 2158
rect 14989 1749 15251 1761
rect 15367 2158 15629 2170
rect 15367 1761 15373 2158
rect 15623 1761 15629 2158
rect 15367 1749 15629 1761
rect 15745 2158 16007 2170
rect 15745 1761 15751 2158
rect 16001 1761 16007 2158
rect 15745 1749 16007 1761
rect 16123 2158 16385 2170
rect 16123 1761 16129 2158
rect 16379 1761 16385 2158
rect 16123 1749 16385 1761
rect 16501 2158 16763 2170
rect 16501 1761 16507 2158
rect 16757 1761 16763 2158
rect 16501 1749 16763 1761
rect 16879 2158 17141 2170
rect 16879 1761 16885 2158
rect 17135 1761 17141 2158
rect 16879 1749 17141 1761
rect 17257 2158 17519 2170
rect 17257 1761 17263 2158
rect 17513 1761 17519 2158
rect 17257 1749 17519 1761
rect 17635 2158 17897 2170
rect 17635 1761 17641 2158
rect 17891 1761 17897 2158
rect 17635 1749 17897 1761
rect 18013 2158 18275 2170
rect 18013 1761 18019 2158
rect 18269 1761 18275 2158
rect 18013 1749 18275 1761
rect 18391 2158 18653 2170
rect 18391 1761 18397 2158
rect 18647 1761 18653 2158
rect 18391 1749 18653 1761
rect 18769 2158 19031 2170
rect 18769 1761 18775 2158
rect 19025 1761 19031 2158
rect 18769 1749 19031 1761
rect 19147 2158 19409 2170
rect 19147 1761 19153 2158
rect 19403 1761 19409 2158
rect 19147 1749 19409 1761
rect 19525 2158 19787 2170
rect 19525 1761 19531 2158
rect 19781 1761 19787 2158
rect 19525 1749 19787 1761
rect -19787 -1761 -19525 -1749
rect -19787 -2158 -19781 -1761
rect -19531 -2158 -19525 -1761
rect -19787 -2170 -19525 -2158
rect -19409 -1761 -19147 -1749
rect -19409 -2158 -19403 -1761
rect -19153 -2158 -19147 -1761
rect -19409 -2170 -19147 -2158
rect -19031 -1761 -18769 -1749
rect -19031 -2158 -19025 -1761
rect -18775 -2158 -18769 -1761
rect -19031 -2170 -18769 -2158
rect -18653 -1761 -18391 -1749
rect -18653 -2158 -18647 -1761
rect -18397 -2158 -18391 -1761
rect -18653 -2170 -18391 -2158
rect -18275 -1761 -18013 -1749
rect -18275 -2158 -18269 -1761
rect -18019 -2158 -18013 -1761
rect -18275 -2170 -18013 -2158
rect -17897 -1761 -17635 -1749
rect -17897 -2158 -17891 -1761
rect -17641 -2158 -17635 -1761
rect -17897 -2170 -17635 -2158
rect -17519 -1761 -17257 -1749
rect -17519 -2158 -17513 -1761
rect -17263 -2158 -17257 -1761
rect -17519 -2170 -17257 -2158
rect -17141 -1761 -16879 -1749
rect -17141 -2158 -17135 -1761
rect -16885 -2158 -16879 -1761
rect -17141 -2170 -16879 -2158
rect -16763 -1761 -16501 -1749
rect -16763 -2158 -16757 -1761
rect -16507 -2158 -16501 -1761
rect -16763 -2170 -16501 -2158
rect -16385 -1761 -16123 -1749
rect -16385 -2158 -16379 -1761
rect -16129 -2158 -16123 -1761
rect -16385 -2170 -16123 -2158
rect -16007 -1761 -15745 -1749
rect -16007 -2158 -16001 -1761
rect -15751 -2158 -15745 -1761
rect -16007 -2170 -15745 -2158
rect -15629 -1761 -15367 -1749
rect -15629 -2158 -15623 -1761
rect -15373 -2158 -15367 -1761
rect -15629 -2170 -15367 -2158
rect -15251 -1761 -14989 -1749
rect -15251 -2158 -15245 -1761
rect -14995 -2158 -14989 -1761
rect -15251 -2170 -14989 -2158
rect -14873 -1761 -14611 -1749
rect -14873 -2158 -14867 -1761
rect -14617 -2158 -14611 -1761
rect -14873 -2170 -14611 -2158
rect -14495 -1761 -14233 -1749
rect -14495 -2158 -14489 -1761
rect -14239 -2158 -14233 -1761
rect -14495 -2170 -14233 -2158
rect -14117 -1761 -13855 -1749
rect -14117 -2158 -14111 -1761
rect -13861 -2158 -13855 -1761
rect -14117 -2170 -13855 -2158
rect -13739 -1761 -13477 -1749
rect -13739 -2158 -13733 -1761
rect -13483 -2158 -13477 -1761
rect -13739 -2170 -13477 -2158
rect -13361 -1761 -13099 -1749
rect -13361 -2158 -13355 -1761
rect -13105 -2158 -13099 -1761
rect -13361 -2170 -13099 -2158
rect -12983 -1761 -12721 -1749
rect -12983 -2158 -12977 -1761
rect -12727 -2158 -12721 -1761
rect -12983 -2170 -12721 -2158
rect -12605 -1761 -12343 -1749
rect -12605 -2158 -12599 -1761
rect -12349 -2158 -12343 -1761
rect -12605 -2170 -12343 -2158
rect -12227 -1761 -11965 -1749
rect -12227 -2158 -12221 -1761
rect -11971 -2158 -11965 -1761
rect -12227 -2170 -11965 -2158
rect -11849 -1761 -11587 -1749
rect -11849 -2158 -11843 -1761
rect -11593 -2158 -11587 -1761
rect -11849 -2170 -11587 -2158
rect -11471 -1761 -11209 -1749
rect -11471 -2158 -11465 -1761
rect -11215 -2158 -11209 -1761
rect -11471 -2170 -11209 -2158
rect -11093 -1761 -10831 -1749
rect -11093 -2158 -11087 -1761
rect -10837 -2158 -10831 -1761
rect -11093 -2170 -10831 -2158
rect -10715 -1761 -10453 -1749
rect -10715 -2158 -10709 -1761
rect -10459 -2158 -10453 -1761
rect -10715 -2170 -10453 -2158
rect -10337 -1761 -10075 -1749
rect -10337 -2158 -10331 -1761
rect -10081 -2158 -10075 -1761
rect -10337 -2170 -10075 -2158
rect -9959 -1761 -9697 -1749
rect -9959 -2158 -9953 -1761
rect -9703 -2158 -9697 -1761
rect -9959 -2170 -9697 -2158
rect -9581 -1761 -9319 -1749
rect -9581 -2158 -9575 -1761
rect -9325 -2158 -9319 -1761
rect -9581 -2170 -9319 -2158
rect -9203 -1761 -8941 -1749
rect -9203 -2158 -9197 -1761
rect -8947 -2158 -8941 -1761
rect -9203 -2170 -8941 -2158
rect -8825 -1761 -8563 -1749
rect -8825 -2158 -8819 -1761
rect -8569 -2158 -8563 -1761
rect -8825 -2170 -8563 -2158
rect -8447 -1761 -8185 -1749
rect -8447 -2158 -8441 -1761
rect -8191 -2158 -8185 -1761
rect -8447 -2170 -8185 -2158
rect -8069 -1761 -7807 -1749
rect -8069 -2158 -8063 -1761
rect -7813 -2158 -7807 -1761
rect -8069 -2170 -7807 -2158
rect -7691 -1761 -7429 -1749
rect -7691 -2158 -7685 -1761
rect -7435 -2158 -7429 -1761
rect -7691 -2170 -7429 -2158
rect -7313 -1761 -7051 -1749
rect -7313 -2158 -7307 -1761
rect -7057 -2158 -7051 -1761
rect -7313 -2170 -7051 -2158
rect -6935 -1761 -6673 -1749
rect -6935 -2158 -6929 -1761
rect -6679 -2158 -6673 -1761
rect -6935 -2170 -6673 -2158
rect -6557 -1761 -6295 -1749
rect -6557 -2158 -6551 -1761
rect -6301 -2158 -6295 -1761
rect -6557 -2170 -6295 -2158
rect -6179 -1761 -5917 -1749
rect -6179 -2158 -6173 -1761
rect -5923 -2158 -5917 -1761
rect -6179 -2170 -5917 -2158
rect -5801 -1761 -5539 -1749
rect -5801 -2158 -5795 -1761
rect -5545 -2158 -5539 -1761
rect -5801 -2170 -5539 -2158
rect -5423 -1761 -5161 -1749
rect -5423 -2158 -5417 -1761
rect -5167 -2158 -5161 -1761
rect -5423 -2170 -5161 -2158
rect -5045 -1761 -4783 -1749
rect -5045 -2158 -5039 -1761
rect -4789 -2158 -4783 -1761
rect -5045 -2170 -4783 -2158
rect -4667 -1761 -4405 -1749
rect -4667 -2158 -4661 -1761
rect -4411 -2158 -4405 -1761
rect -4667 -2170 -4405 -2158
rect -4289 -1761 -4027 -1749
rect -4289 -2158 -4283 -1761
rect -4033 -2158 -4027 -1761
rect -4289 -2170 -4027 -2158
rect -3911 -1761 -3649 -1749
rect -3911 -2158 -3905 -1761
rect -3655 -2158 -3649 -1761
rect -3911 -2170 -3649 -2158
rect -3533 -1761 -3271 -1749
rect -3533 -2158 -3527 -1761
rect -3277 -2158 -3271 -1761
rect -3533 -2170 -3271 -2158
rect -3155 -1761 -2893 -1749
rect -3155 -2158 -3149 -1761
rect -2899 -2158 -2893 -1761
rect -3155 -2170 -2893 -2158
rect -2777 -1761 -2515 -1749
rect -2777 -2158 -2771 -1761
rect -2521 -2158 -2515 -1761
rect -2777 -2170 -2515 -2158
rect -2399 -1761 -2137 -1749
rect -2399 -2158 -2393 -1761
rect -2143 -2158 -2137 -1761
rect -2399 -2170 -2137 -2158
rect -2021 -1761 -1759 -1749
rect -2021 -2158 -2015 -1761
rect -1765 -2158 -1759 -1761
rect -2021 -2170 -1759 -2158
rect -1643 -1761 -1381 -1749
rect -1643 -2158 -1637 -1761
rect -1387 -2158 -1381 -1761
rect -1643 -2170 -1381 -2158
rect -1265 -1761 -1003 -1749
rect -1265 -2158 -1259 -1761
rect -1009 -2158 -1003 -1761
rect -1265 -2170 -1003 -2158
rect -887 -1761 -625 -1749
rect -887 -2158 -881 -1761
rect -631 -2158 -625 -1761
rect -887 -2170 -625 -2158
rect -509 -1761 -247 -1749
rect -509 -2158 -503 -1761
rect -253 -2158 -247 -1761
rect -509 -2170 -247 -2158
rect -131 -1761 131 -1749
rect -131 -2158 -125 -1761
rect 125 -2158 131 -1761
rect -131 -2170 131 -2158
rect 247 -1761 509 -1749
rect 247 -2158 253 -1761
rect 503 -2158 509 -1761
rect 247 -2170 509 -2158
rect 625 -1761 887 -1749
rect 625 -2158 631 -1761
rect 881 -2158 887 -1761
rect 625 -2170 887 -2158
rect 1003 -1761 1265 -1749
rect 1003 -2158 1009 -1761
rect 1259 -2158 1265 -1761
rect 1003 -2170 1265 -2158
rect 1381 -1761 1643 -1749
rect 1381 -2158 1387 -1761
rect 1637 -2158 1643 -1761
rect 1381 -2170 1643 -2158
rect 1759 -1761 2021 -1749
rect 1759 -2158 1765 -1761
rect 2015 -2158 2021 -1761
rect 1759 -2170 2021 -2158
rect 2137 -1761 2399 -1749
rect 2137 -2158 2143 -1761
rect 2393 -2158 2399 -1761
rect 2137 -2170 2399 -2158
rect 2515 -1761 2777 -1749
rect 2515 -2158 2521 -1761
rect 2771 -2158 2777 -1761
rect 2515 -2170 2777 -2158
rect 2893 -1761 3155 -1749
rect 2893 -2158 2899 -1761
rect 3149 -2158 3155 -1761
rect 2893 -2170 3155 -2158
rect 3271 -1761 3533 -1749
rect 3271 -2158 3277 -1761
rect 3527 -2158 3533 -1761
rect 3271 -2170 3533 -2158
rect 3649 -1761 3911 -1749
rect 3649 -2158 3655 -1761
rect 3905 -2158 3911 -1761
rect 3649 -2170 3911 -2158
rect 4027 -1761 4289 -1749
rect 4027 -2158 4033 -1761
rect 4283 -2158 4289 -1761
rect 4027 -2170 4289 -2158
rect 4405 -1761 4667 -1749
rect 4405 -2158 4411 -1761
rect 4661 -2158 4667 -1761
rect 4405 -2170 4667 -2158
rect 4783 -1761 5045 -1749
rect 4783 -2158 4789 -1761
rect 5039 -2158 5045 -1761
rect 4783 -2170 5045 -2158
rect 5161 -1761 5423 -1749
rect 5161 -2158 5167 -1761
rect 5417 -2158 5423 -1761
rect 5161 -2170 5423 -2158
rect 5539 -1761 5801 -1749
rect 5539 -2158 5545 -1761
rect 5795 -2158 5801 -1761
rect 5539 -2170 5801 -2158
rect 5917 -1761 6179 -1749
rect 5917 -2158 5923 -1761
rect 6173 -2158 6179 -1761
rect 5917 -2170 6179 -2158
rect 6295 -1761 6557 -1749
rect 6295 -2158 6301 -1761
rect 6551 -2158 6557 -1761
rect 6295 -2170 6557 -2158
rect 6673 -1761 6935 -1749
rect 6673 -2158 6679 -1761
rect 6929 -2158 6935 -1761
rect 6673 -2170 6935 -2158
rect 7051 -1761 7313 -1749
rect 7051 -2158 7057 -1761
rect 7307 -2158 7313 -1761
rect 7051 -2170 7313 -2158
rect 7429 -1761 7691 -1749
rect 7429 -2158 7435 -1761
rect 7685 -2158 7691 -1761
rect 7429 -2170 7691 -2158
rect 7807 -1761 8069 -1749
rect 7807 -2158 7813 -1761
rect 8063 -2158 8069 -1761
rect 7807 -2170 8069 -2158
rect 8185 -1761 8447 -1749
rect 8185 -2158 8191 -1761
rect 8441 -2158 8447 -1761
rect 8185 -2170 8447 -2158
rect 8563 -1761 8825 -1749
rect 8563 -2158 8569 -1761
rect 8819 -2158 8825 -1761
rect 8563 -2170 8825 -2158
rect 8941 -1761 9203 -1749
rect 8941 -2158 8947 -1761
rect 9197 -2158 9203 -1761
rect 8941 -2170 9203 -2158
rect 9319 -1761 9581 -1749
rect 9319 -2158 9325 -1761
rect 9575 -2158 9581 -1761
rect 9319 -2170 9581 -2158
rect 9697 -1761 9959 -1749
rect 9697 -2158 9703 -1761
rect 9953 -2158 9959 -1761
rect 9697 -2170 9959 -2158
rect 10075 -1761 10337 -1749
rect 10075 -2158 10081 -1761
rect 10331 -2158 10337 -1761
rect 10075 -2170 10337 -2158
rect 10453 -1761 10715 -1749
rect 10453 -2158 10459 -1761
rect 10709 -2158 10715 -1761
rect 10453 -2170 10715 -2158
rect 10831 -1761 11093 -1749
rect 10831 -2158 10837 -1761
rect 11087 -2158 11093 -1761
rect 10831 -2170 11093 -2158
rect 11209 -1761 11471 -1749
rect 11209 -2158 11215 -1761
rect 11465 -2158 11471 -1761
rect 11209 -2170 11471 -2158
rect 11587 -1761 11849 -1749
rect 11587 -2158 11593 -1761
rect 11843 -2158 11849 -1761
rect 11587 -2170 11849 -2158
rect 11965 -1761 12227 -1749
rect 11965 -2158 11971 -1761
rect 12221 -2158 12227 -1761
rect 11965 -2170 12227 -2158
rect 12343 -1761 12605 -1749
rect 12343 -2158 12349 -1761
rect 12599 -2158 12605 -1761
rect 12343 -2170 12605 -2158
rect 12721 -1761 12983 -1749
rect 12721 -2158 12727 -1761
rect 12977 -2158 12983 -1761
rect 12721 -2170 12983 -2158
rect 13099 -1761 13361 -1749
rect 13099 -2158 13105 -1761
rect 13355 -2158 13361 -1761
rect 13099 -2170 13361 -2158
rect 13477 -1761 13739 -1749
rect 13477 -2158 13483 -1761
rect 13733 -2158 13739 -1761
rect 13477 -2170 13739 -2158
rect 13855 -1761 14117 -1749
rect 13855 -2158 13861 -1761
rect 14111 -2158 14117 -1761
rect 13855 -2170 14117 -2158
rect 14233 -1761 14495 -1749
rect 14233 -2158 14239 -1761
rect 14489 -2158 14495 -1761
rect 14233 -2170 14495 -2158
rect 14611 -1761 14873 -1749
rect 14611 -2158 14617 -1761
rect 14867 -2158 14873 -1761
rect 14611 -2170 14873 -2158
rect 14989 -1761 15251 -1749
rect 14989 -2158 14995 -1761
rect 15245 -2158 15251 -1761
rect 14989 -2170 15251 -2158
rect 15367 -1761 15629 -1749
rect 15367 -2158 15373 -1761
rect 15623 -2158 15629 -1761
rect 15367 -2170 15629 -2158
rect 15745 -1761 16007 -1749
rect 15745 -2158 15751 -1761
rect 16001 -2158 16007 -1761
rect 15745 -2170 16007 -2158
rect 16123 -1761 16385 -1749
rect 16123 -2158 16129 -1761
rect 16379 -2158 16385 -1761
rect 16123 -2170 16385 -2158
rect 16501 -1761 16763 -1749
rect 16501 -2158 16507 -1761
rect 16757 -2158 16763 -1761
rect 16501 -2170 16763 -2158
rect 16879 -1761 17141 -1749
rect 16879 -2158 16885 -1761
rect 17135 -2158 17141 -1761
rect 16879 -2170 17141 -2158
rect 17257 -1761 17519 -1749
rect 17257 -2158 17263 -1761
rect 17513 -2158 17519 -1761
rect 17257 -2170 17519 -2158
rect 17635 -1761 17897 -1749
rect 17635 -2158 17641 -1761
rect 17891 -2158 17897 -1761
rect 17635 -2170 17897 -2158
rect 18013 -1761 18275 -1749
rect 18013 -2158 18019 -1761
rect 18269 -2158 18275 -1761
rect 18013 -2170 18275 -2158
rect 18391 -1761 18653 -1749
rect 18391 -2158 18397 -1761
rect 18647 -2158 18653 -1761
rect 18391 -2170 18653 -2158
rect 18769 -1761 19031 -1749
rect 18769 -2158 18775 -1761
rect 19025 -2158 19031 -1761
rect 18769 -2170 19031 -2158
rect 19147 -1761 19409 -1749
rect 19147 -2158 19153 -1761
rect 19403 -2158 19409 -1761
rect 19147 -2170 19409 -2158
rect 19525 -1761 19787 -1749
rect 19525 -2158 19531 -1761
rect 19781 -2158 19787 -1761
rect 19525 -2170 19787 -2158
<< properties >>
string FIXED_BBOX -19931 -2310 19931 2310
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.41 l 17.6 m 1 nx 105 wmin 1.410 lmin 0.50 rho 2000 val 25.231k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 1 hv_guard 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
