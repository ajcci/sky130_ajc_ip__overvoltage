magic
tech sky130A
magscale 1 2
timestamp 1711600228
<< mvnmos >>
rect -60 -531 60 469
<< mvndiff >>
rect -118 457 -60 469
rect -118 -519 -106 457
rect -72 -519 -60 457
rect -118 -531 -60 -519
rect 60 457 118 469
rect 60 -519 72 457
rect 106 -519 118 457
rect 60 -531 118 -519
<< mvndiffc >>
rect -106 -519 -72 457
rect 72 -519 106 457
<< poly >>
rect -60 541 60 557
rect -60 507 -44 541
rect 44 507 60 541
rect -60 469 60 507
rect -60 -557 60 -531
<< polycont >>
rect -44 507 44 541
<< locali >>
rect -60 507 -44 541
rect 44 507 60 541
rect -106 457 -72 473
rect -106 -535 -72 -519
rect 72 457 106 473
rect 72 -535 106 -519
<< viali >>
rect -44 507 44 541
rect -106 -519 -72 457
rect 72 -519 106 457
<< metal1 >>
rect -56 541 56 547
rect -56 507 -44 541
rect 44 507 56 541
rect -56 501 56 507
rect -112 457 -66 469
rect -112 -519 -106 457
rect -72 -519 -66 457
rect -112 -531 -66 -519
rect 66 457 112 469
rect 66 -519 72 457
rect 106 -519 112 457
rect 66 -531 112 -519
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.60 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
