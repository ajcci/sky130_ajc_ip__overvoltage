* SPICE3 file created from comparator.ext - technology: sky130A

*.subckt comparator avdd ibias out ena vinn vinp avss
X0 vt vinn vnn vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X1 vt vinp vpp vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X2 vt vinp vpp vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X3 vt vinp vpp vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X5 vt vinn vnn vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X6 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X7 vt vinp vpp vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X9 vt vinn vnn vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X11 vt vinn vnn vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X12 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X13 vt vinn vnn vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X15 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X16 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X17 vt vinn vnn vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X19 vt vinn vnn vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X20 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X21 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X23 vt vinn vnn vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X24 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X31 vt vinp vpp vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X33 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X34 vt vinp vpp vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X36 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X37 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X38 vt vinp vpp vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X39 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X40 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X41 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X43 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X44 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X46 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X47 vt vinp vpp vt sky130_fd_pr__nfet_g5v0d10v5 w=4.2e-07 l=8e-06
X48 n0 vm avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=8e-06
X49 vm vm avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=8e-06
X51 vt vn avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=8e-06
X53 avss vn vt avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=8e-06
X54 vn vn avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=8e-06
X56 avss vm vm avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=8e-06
X58 avss vm n0 avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=8e-06
X59 avss vn vn avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=8e-06
X60 avdd vnn vm avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=8e-06
X62 n0 vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=8e-06
X63 avdd vpp n0 avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=8e-06
X65 vm vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=8e-06
X66 vnn ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=1e-06
X67 vpp ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=1e-06
X68 ena_b ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=1e-06
X69 vn ena_b ibias avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=1e-06
X70 vn ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=1e-06
X71 vn ena ibias avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=1e-06
X72 n0 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=1e-06
X73 ena_b ena avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=1e-06
X74 vm ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=1e-06
X75 avss n1 out avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X76 avss n1 out avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X77 out n1 avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X78 out n1 avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X79 avss n1 out avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X80 avss n0 n1 avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X81 avss n1 out avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X82 out n1 avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X83 n1 n0 avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X84 out n1 avss avss sky130_fd_pr__nfet_g5v0d10v5 w=1e-06 l=6e-07
X85 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X87 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X91 vnn vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X92 vpp vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X93 vnn vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X94 avdd vpp vnn avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X95 avdd vnn vnn avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X96 avdd vnn vnn avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X97 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X99 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X103 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X104 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X105 avdd vpp vpp avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X108 vpp vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X110 avdd vpp vnn avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X111 avdd vpp vnn avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X113 avdd vnn vpp avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X114 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X115 avdd vnn vpp avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X116 avdd vpp vnn avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X117 avdd vpp vpp avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X118 vpp vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X119 vpp vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X120 vnn vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X121 avdd vnn vpp avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X123 avdd vnn vnn avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X124 avdd vnn vpp avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X127 avdd vpp vpp avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X128 avdd vpp vpp avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X129 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X130 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X132 vnn vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X133 avdd vpp vnn avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X135 avdd vnn vnn avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X137 avdd vnn vpp avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X138 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=4.2e-07 l=8e-06
X139 avdd n0 n1 avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
X140 avdd n1 out avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
X141 out n1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
X142 n1 n0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
X143 out n1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
X144 avdd n1 out avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
X145 avdd n1 out avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
X146 out n1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
X147 out n1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
X148 avdd n1 out avdd sky130_fd_pr__pfet_g5v0d10v5 w=1e-06 l=6e-07
*.ends
