magic
tech sky130A
magscale 1 2
timestamp 1712337786
<< error_s >>
rect 41712 -6012 42971 -6011
rect 41712 -6015 42976 -6012
rect 41703 -6016 42976 -6015
rect 41698 -6054 42976 -6016
rect 41694 -6063 41776 -6054
rect 42906 -6063 42911 -6054
rect 42915 -6059 42971 -6054
rect 42975 -6063 42980 -6054
rect 41703 -6080 41767 -6063
rect 47737 -6108 47802 -6049
rect 47736 -6109 47802 -6108
rect 47736 -6113 47797 -6109
rect 47736 -6169 47741 -6113
rect 47792 -6114 47797 -6113
rect 47792 -6169 47802 -6114
rect 47736 -6174 47802 -6169
rect 48265 -6292 48330 -6233
rect 48264 -6293 48330 -6292
rect 48264 -6297 48325 -6293
rect 48264 -6353 48269 -6297
rect 48320 -6298 48325 -6297
rect 48320 -6353 48330 -6298
rect 48264 -6358 48330 -6353
rect 48795 -6439 48860 -6380
rect 48794 -6440 48860 -6439
rect 48794 -6444 48855 -6440
rect 48794 -6500 48799 -6444
rect 48850 -6445 48855 -6444
rect 48850 -6500 48860 -6445
rect 48794 -6505 48860 -6500
<< metal1 >>
rect 35387 -10127 40107 -10121
rect 35387 -10315 39918 -10127
rect 40101 -10315 40107 -10127
rect 35387 -10321 40107 -10315
rect 35387 -10577 40357 -10377
<< via1 >>
rect 40420 -6997 40608 -6861
rect 39918 -10315 40101 -10127
rect 40419 -10315 40607 -10127
<< metal2 >>
rect 40414 -6861 40614 -6054
rect 41703 -6080 41767 -6071
rect 42911 -6067 42915 -6054
rect 42971 -6067 42975 -6054
rect 42380 -6173 42436 -6168
rect 42376 -6177 42440 -6173
rect 42376 -6233 42380 -6177
rect 42436 -6233 42440 -6177
rect 41852 -6311 41908 -6306
rect 41848 -6315 41912 -6311
rect 41848 -6371 41852 -6315
rect 41908 -6371 41912 -6315
rect 41328 -6449 41384 -6444
rect 41324 -6453 41388 -6449
rect 41324 -6509 41328 -6453
rect 41384 -6509 41388 -6453
rect 40782 -6599 40838 -6590
rect 40782 -6664 40838 -6655
rect 41324 -6668 41388 -6509
rect 41848 -6679 41912 -6371
rect 42376 -6671 42440 -6233
rect 42911 -6671 42975 -6067
rect 43461 -6671 43525 -6054
rect 43815 -6600 43879 -6054
rect 43974 -6419 44038 -6054
rect 44528 -6419 44584 -6414
rect 43974 -6492 44038 -6483
rect 44524 -6423 44588 -6419
rect 44524 -6479 44528 -6423
rect 44584 -6479 44588 -6423
rect 43815 -6664 44060 -6600
rect 44524 -6679 44588 -6479
rect 45066 -6671 45130 -6061
rect 45587 -6664 45651 -6061
rect 46130 -6629 46194 -6061
rect 46659 -6672 46723 -6061
rect 47195 -6679 47259 -6061
rect 47741 -6109 47797 -6104
rect 47737 -6113 47801 -6109
rect 47737 -6169 47741 -6113
rect 47797 -6169 47801 -6113
rect 47737 -6687 47801 -6169
rect 48269 -6293 48325 -6288
rect 48265 -6297 48329 -6293
rect 48265 -6353 48269 -6297
rect 48325 -6353 48329 -6297
rect 48265 -6665 48329 -6353
rect 48799 -6440 48855 -6435
rect 48795 -6444 48859 -6440
rect 48795 -6500 48799 -6444
rect 48855 -6500 48859 -6444
rect 48795 -6665 48859 -6500
rect 48955 -6687 49019 -6545
rect 40414 -6997 40420 -6861
rect 40608 -6997 40614 -6861
rect 40414 -7003 40614 -6997
rect 40604 -7339 40664 -7330
rect 39906 -8077 39970 -7555
rect 40604 -8201 40664 -7399
rect 40604 -8257 40606 -8201
rect 40662 -8257 40664 -8201
rect 40604 -8259 40664 -8257
rect 40606 -8266 40662 -8259
rect 39912 -10127 40613 -10121
rect 39912 -10315 39918 -10127
rect 40101 -10315 40419 -10127
rect 40607 -10315 40613 -10127
rect 39912 -10321 40613 -10315
<< via2 >>
rect 41703 -6071 41767 -6054
rect 42915 -6067 42971 -6054
rect 42380 -6233 42436 -6177
rect 41852 -6371 41908 -6315
rect 41328 -6509 41384 -6453
rect 40782 -6655 40838 -6599
rect 43974 -6483 44038 -6419
rect 44528 -6479 44584 -6423
rect 47741 -6169 47797 -6113
rect 48269 -6353 48325 -6297
rect 48799 -6500 48855 -6444
rect 40604 -7399 40664 -7339
rect 40606 -8257 40662 -8201
<< metal3 >>
rect 41698 -6071 41703 -6054
rect 41767 -6067 42915 -6054
rect 42971 -6067 42976 -6054
rect 41767 -6071 42976 -6067
rect 41698 -6076 41772 -6071
rect 42910 -6072 42976 -6071
rect 47736 -6109 47802 -6108
rect 47736 -6113 47797 -6109
rect 47736 -6169 47741 -6113
rect 42375 -6173 42441 -6172
rect 40151 -6177 42441 -6173
rect 47736 -6173 47797 -6169
rect 47736 -6174 47802 -6173
rect 40151 -6233 42380 -6177
rect 42436 -6233 42441 -6177
rect 40151 -6237 42441 -6233
rect 42375 -6238 42441 -6237
rect 48264 -6293 48330 -6292
rect 48264 -6297 48325 -6293
rect 41847 -6311 41913 -6310
rect 40151 -6315 41913 -6311
rect 40151 -6371 41852 -6315
rect 41908 -6371 41913 -6315
rect 48264 -6353 48269 -6297
rect 48264 -6357 48325 -6353
rect 48264 -6358 48330 -6357
rect 40151 -6375 41913 -6371
rect 41847 -6376 41913 -6375
rect 43969 -6419 44043 -6414
rect 44523 -6419 44589 -6418
rect 41323 -6449 41389 -6448
rect 40151 -6453 41389 -6449
rect 40151 -6509 41328 -6453
rect 41384 -6509 41389 -6453
rect 43969 -6483 43974 -6419
rect 44038 -6423 44589 -6419
rect 44038 -6479 44528 -6423
rect 44584 -6479 44589 -6423
rect 44038 -6483 44589 -6479
rect 43969 -6488 44043 -6483
rect 44523 -6484 44589 -6483
rect 48794 -6440 48860 -6439
rect 48794 -6444 48855 -6440
rect 48794 -6500 48799 -6444
rect 48794 -6504 48855 -6500
rect 48794 -6505 48860 -6504
rect 40151 -6513 41389 -6509
rect 41323 -6514 41389 -6513
rect 40777 -6595 40843 -6594
rect 40151 -6599 40843 -6595
rect 40151 -6655 40782 -6599
rect 40838 -6655 40843 -6599
rect 40151 -6659 40843 -6655
rect 40777 -6660 40843 -6659
rect 40599 -7339 40669 -7334
rect 40151 -7399 40604 -7339
rect 40664 -7399 40669 -7339
rect 40599 -7404 40669 -7399
rect 40601 -8199 40667 -8196
rect 40601 -8201 41265 -8199
rect 40601 -8257 40606 -8201
rect 40662 -8257 41265 -8201
rect 40601 -8259 41265 -8257
rect 48718 -8259 48778 -8199
rect 40601 -8262 40667 -8259
use rstring_mux  rstring_mux_0
timestamp 1712334093
transform 1 0 28241 0 1 -15265
box -11632 -32 28451 9182
<< end >>
