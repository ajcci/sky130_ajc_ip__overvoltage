xspice/overvoltage_dig.out.spice