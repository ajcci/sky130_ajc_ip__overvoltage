magic
tech sky130A
magscale 1 2
timestamp 1712158818
<< pwell >>
rect -4382 -727 4382 727
<< mvnmos >>
rect -4154 -469 -4034 531
rect -3976 -469 -3856 531
rect -3798 -469 -3678 531
rect -3620 -469 -3500 531
rect -3442 -469 -3322 531
rect -3264 -469 -3144 531
rect -3086 -469 -2966 531
rect -2908 -469 -2788 531
rect -2730 -469 -2610 531
rect -2552 -469 -2432 531
rect -2374 -469 -2254 531
rect -2196 -469 -2076 531
rect -2018 -469 -1898 531
rect -1840 -469 -1720 531
rect -1662 -469 -1542 531
rect -1484 -469 -1364 531
rect -1306 -469 -1186 531
rect -1128 -469 -1008 531
rect -950 -469 -830 531
rect -772 -469 -652 531
rect -594 -469 -474 531
rect -416 -469 -296 531
rect -238 -469 -118 531
rect -60 -469 60 531
rect 118 -469 238 531
rect 296 -469 416 531
rect 474 -469 594 531
rect 652 -469 772 531
rect 830 -469 950 531
rect 1008 -469 1128 531
rect 1186 -469 1306 531
rect 1364 -469 1484 531
rect 1542 -469 1662 531
rect 1720 -469 1840 531
rect 1898 -469 2018 531
rect 2076 -469 2196 531
rect 2254 -469 2374 531
rect 2432 -469 2552 531
rect 2610 -469 2730 531
rect 2788 -469 2908 531
rect 2966 -469 3086 531
rect 3144 -469 3264 531
rect 3322 -469 3442 531
rect 3500 -469 3620 531
rect 3678 -469 3798 531
rect 3856 -469 3976 531
rect 4034 -469 4154 531
<< mvndiff >>
rect -4212 519 -4154 531
rect -4212 -457 -4200 519
rect -4166 -457 -4154 519
rect -4212 -469 -4154 -457
rect -4034 519 -3976 531
rect -4034 -457 -4022 519
rect -3988 -457 -3976 519
rect -4034 -469 -3976 -457
rect -3856 519 -3798 531
rect -3856 -457 -3844 519
rect -3810 -457 -3798 519
rect -3856 -469 -3798 -457
rect -3678 519 -3620 531
rect -3678 -457 -3666 519
rect -3632 -457 -3620 519
rect -3678 -469 -3620 -457
rect -3500 519 -3442 531
rect -3500 -457 -3488 519
rect -3454 -457 -3442 519
rect -3500 -469 -3442 -457
rect -3322 519 -3264 531
rect -3322 -457 -3310 519
rect -3276 -457 -3264 519
rect -3322 -469 -3264 -457
rect -3144 519 -3086 531
rect -3144 -457 -3132 519
rect -3098 -457 -3086 519
rect -3144 -469 -3086 -457
rect -2966 519 -2908 531
rect -2966 -457 -2954 519
rect -2920 -457 -2908 519
rect -2966 -469 -2908 -457
rect -2788 519 -2730 531
rect -2788 -457 -2776 519
rect -2742 -457 -2730 519
rect -2788 -469 -2730 -457
rect -2610 519 -2552 531
rect -2610 -457 -2598 519
rect -2564 -457 -2552 519
rect -2610 -469 -2552 -457
rect -2432 519 -2374 531
rect -2432 -457 -2420 519
rect -2386 -457 -2374 519
rect -2432 -469 -2374 -457
rect -2254 519 -2196 531
rect -2254 -457 -2242 519
rect -2208 -457 -2196 519
rect -2254 -469 -2196 -457
rect -2076 519 -2018 531
rect -2076 -457 -2064 519
rect -2030 -457 -2018 519
rect -2076 -469 -2018 -457
rect -1898 519 -1840 531
rect -1898 -457 -1886 519
rect -1852 -457 -1840 519
rect -1898 -469 -1840 -457
rect -1720 519 -1662 531
rect -1720 -457 -1708 519
rect -1674 -457 -1662 519
rect -1720 -469 -1662 -457
rect -1542 519 -1484 531
rect -1542 -457 -1530 519
rect -1496 -457 -1484 519
rect -1542 -469 -1484 -457
rect -1364 519 -1306 531
rect -1364 -457 -1352 519
rect -1318 -457 -1306 519
rect -1364 -469 -1306 -457
rect -1186 519 -1128 531
rect -1186 -457 -1174 519
rect -1140 -457 -1128 519
rect -1186 -469 -1128 -457
rect -1008 519 -950 531
rect -1008 -457 -996 519
rect -962 -457 -950 519
rect -1008 -469 -950 -457
rect -830 519 -772 531
rect -830 -457 -818 519
rect -784 -457 -772 519
rect -830 -469 -772 -457
rect -652 519 -594 531
rect -652 -457 -640 519
rect -606 -457 -594 519
rect -652 -469 -594 -457
rect -474 519 -416 531
rect -474 -457 -462 519
rect -428 -457 -416 519
rect -474 -469 -416 -457
rect -296 519 -238 531
rect -296 -457 -284 519
rect -250 -457 -238 519
rect -296 -469 -238 -457
rect -118 519 -60 531
rect -118 -457 -106 519
rect -72 -457 -60 519
rect -118 -469 -60 -457
rect 60 519 118 531
rect 60 -457 72 519
rect 106 -457 118 519
rect 60 -469 118 -457
rect 238 519 296 531
rect 238 -457 250 519
rect 284 -457 296 519
rect 238 -469 296 -457
rect 416 519 474 531
rect 416 -457 428 519
rect 462 -457 474 519
rect 416 -469 474 -457
rect 594 519 652 531
rect 594 -457 606 519
rect 640 -457 652 519
rect 594 -469 652 -457
rect 772 519 830 531
rect 772 -457 784 519
rect 818 -457 830 519
rect 772 -469 830 -457
rect 950 519 1008 531
rect 950 -457 962 519
rect 996 -457 1008 519
rect 950 -469 1008 -457
rect 1128 519 1186 531
rect 1128 -457 1140 519
rect 1174 -457 1186 519
rect 1128 -469 1186 -457
rect 1306 519 1364 531
rect 1306 -457 1318 519
rect 1352 -457 1364 519
rect 1306 -469 1364 -457
rect 1484 519 1542 531
rect 1484 -457 1496 519
rect 1530 -457 1542 519
rect 1484 -469 1542 -457
rect 1662 519 1720 531
rect 1662 -457 1674 519
rect 1708 -457 1720 519
rect 1662 -469 1720 -457
rect 1840 519 1898 531
rect 1840 -457 1852 519
rect 1886 -457 1898 519
rect 1840 -469 1898 -457
rect 2018 519 2076 531
rect 2018 -457 2030 519
rect 2064 -457 2076 519
rect 2018 -469 2076 -457
rect 2196 519 2254 531
rect 2196 -457 2208 519
rect 2242 -457 2254 519
rect 2196 -469 2254 -457
rect 2374 519 2432 531
rect 2374 -457 2386 519
rect 2420 -457 2432 519
rect 2374 -469 2432 -457
rect 2552 519 2610 531
rect 2552 -457 2564 519
rect 2598 -457 2610 519
rect 2552 -469 2610 -457
rect 2730 519 2788 531
rect 2730 -457 2742 519
rect 2776 -457 2788 519
rect 2730 -469 2788 -457
rect 2908 519 2966 531
rect 2908 -457 2920 519
rect 2954 -457 2966 519
rect 2908 -469 2966 -457
rect 3086 519 3144 531
rect 3086 -457 3098 519
rect 3132 -457 3144 519
rect 3086 -469 3144 -457
rect 3264 519 3322 531
rect 3264 -457 3276 519
rect 3310 -457 3322 519
rect 3264 -469 3322 -457
rect 3442 519 3500 531
rect 3442 -457 3454 519
rect 3488 -457 3500 519
rect 3442 -469 3500 -457
rect 3620 519 3678 531
rect 3620 -457 3632 519
rect 3666 -457 3678 519
rect 3620 -469 3678 -457
rect 3798 519 3856 531
rect 3798 -457 3810 519
rect 3844 -457 3856 519
rect 3798 -469 3856 -457
rect 3976 519 4034 531
rect 3976 -457 3988 519
rect 4022 -457 4034 519
rect 3976 -469 4034 -457
rect 4154 519 4212 531
rect 4154 -457 4166 519
rect 4200 -457 4212 519
rect 4154 -469 4212 -457
<< mvndiffc >>
rect -4200 -457 -4166 519
rect -4022 -457 -3988 519
rect -3844 -457 -3810 519
rect -3666 -457 -3632 519
rect -3488 -457 -3454 519
rect -3310 -457 -3276 519
rect -3132 -457 -3098 519
rect -2954 -457 -2920 519
rect -2776 -457 -2742 519
rect -2598 -457 -2564 519
rect -2420 -457 -2386 519
rect -2242 -457 -2208 519
rect -2064 -457 -2030 519
rect -1886 -457 -1852 519
rect -1708 -457 -1674 519
rect -1530 -457 -1496 519
rect -1352 -457 -1318 519
rect -1174 -457 -1140 519
rect -996 -457 -962 519
rect -818 -457 -784 519
rect -640 -457 -606 519
rect -462 -457 -428 519
rect -284 -457 -250 519
rect -106 -457 -72 519
rect 72 -457 106 519
rect 250 -457 284 519
rect 428 -457 462 519
rect 606 -457 640 519
rect 784 -457 818 519
rect 962 -457 996 519
rect 1140 -457 1174 519
rect 1318 -457 1352 519
rect 1496 -457 1530 519
rect 1674 -457 1708 519
rect 1852 -457 1886 519
rect 2030 -457 2064 519
rect 2208 -457 2242 519
rect 2386 -457 2420 519
rect 2564 -457 2598 519
rect 2742 -457 2776 519
rect 2920 -457 2954 519
rect 3098 -457 3132 519
rect 3276 -457 3310 519
rect 3454 -457 3488 519
rect 3632 -457 3666 519
rect 3810 -457 3844 519
rect 3988 -457 4022 519
rect 4166 -457 4200 519
<< mvpsubdiff >>
rect -4346 679 4346 691
rect -4346 645 -4238 679
rect 4238 645 4346 679
rect -4346 633 4346 645
rect -4346 583 -4288 633
rect -4346 -583 -4334 583
rect -4300 -583 -4288 583
rect 4288 583 4346 633
rect -4346 -633 -4288 -583
rect 4288 -583 4300 583
rect 4334 -583 4346 583
rect 4288 -633 4346 -583
rect -4346 -645 4346 -633
rect -4346 -679 -4238 -645
rect 4238 -679 4346 -645
rect -4346 -691 4346 -679
<< mvpsubdiffcont >>
rect -4238 645 4238 679
rect -4334 -583 -4300 583
rect 4300 -583 4334 583
rect -4238 -679 4238 -645
<< poly >>
rect -4154 531 -4034 557
rect -3976 531 -3856 557
rect -3798 531 -3678 557
rect -3620 531 -3500 557
rect -3442 531 -3322 557
rect -3264 531 -3144 557
rect -3086 531 -2966 557
rect -2908 531 -2788 557
rect -2730 531 -2610 557
rect -2552 531 -2432 557
rect -2374 531 -2254 557
rect -2196 531 -2076 557
rect -2018 531 -1898 557
rect -1840 531 -1720 557
rect -1662 531 -1542 557
rect -1484 531 -1364 557
rect -1306 531 -1186 557
rect -1128 531 -1008 557
rect -950 531 -830 557
rect -772 531 -652 557
rect -594 531 -474 557
rect -416 531 -296 557
rect -238 531 -118 557
rect -60 531 60 557
rect 118 531 238 557
rect 296 531 416 557
rect 474 531 594 557
rect 652 531 772 557
rect 830 531 950 557
rect 1008 531 1128 557
rect 1186 531 1306 557
rect 1364 531 1484 557
rect 1542 531 1662 557
rect 1720 531 1840 557
rect 1898 531 2018 557
rect 2076 531 2196 557
rect 2254 531 2374 557
rect 2432 531 2552 557
rect 2610 531 2730 557
rect 2788 531 2908 557
rect 2966 531 3086 557
rect 3144 531 3264 557
rect 3322 531 3442 557
rect 3500 531 3620 557
rect 3678 531 3798 557
rect 3856 531 3976 557
rect 4034 531 4154 557
rect -4154 -507 -4034 -469
rect -4154 -541 -4138 -507
rect -4050 -541 -4034 -507
rect -4154 -557 -4034 -541
rect -3976 -507 -3856 -469
rect -3976 -541 -3960 -507
rect -3872 -541 -3856 -507
rect -3976 -557 -3856 -541
rect -3798 -507 -3678 -469
rect -3798 -541 -3782 -507
rect -3694 -541 -3678 -507
rect -3798 -557 -3678 -541
rect -3620 -507 -3500 -469
rect -3620 -541 -3604 -507
rect -3516 -541 -3500 -507
rect -3620 -557 -3500 -541
rect -3442 -507 -3322 -469
rect -3442 -541 -3426 -507
rect -3338 -541 -3322 -507
rect -3442 -557 -3322 -541
rect -3264 -507 -3144 -469
rect -3264 -541 -3248 -507
rect -3160 -541 -3144 -507
rect -3264 -557 -3144 -541
rect -3086 -507 -2966 -469
rect -3086 -541 -3070 -507
rect -2982 -541 -2966 -507
rect -3086 -557 -2966 -541
rect -2908 -507 -2788 -469
rect -2908 -541 -2892 -507
rect -2804 -541 -2788 -507
rect -2908 -557 -2788 -541
rect -2730 -507 -2610 -469
rect -2730 -541 -2714 -507
rect -2626 -541 -2610 -507
rect -2730 -557 -2610 -541
rect -2552 -507 -2432 -469
rect -2552 -541 -2536 -507
rect -2448 -541 -2432 -507
rect -2552 -557 -2432 -541
rect -2374 -507 -2254 -469
rect -2374 -541 -2358 -507
rect -2270 -541 -2254 -507
rect -2374 -557 -2254 -541
rect -2196 -507 -2076 -469
rect -2196 -541 -2180 -507
rect -2092 -541 -2076 -507
rect -2196 -557 -2076 -541
rect -2018 -507 -1898 -469
rect -2018 -541 -2002 -507
rect -1914 -541 -1898 -507
rect -2018 -557 -1898 -541
rect -1840 -507 -1720 -469
rect -1840 -541 -1824 -507
rect -1736 -541 -1720 -507
rect -1840 -557 -1720 -541
rect -1662 -507 -1542 -469
rect -1662 -541 -1646 -507
rect -1558 -541 -1542 -507
rect -1662 -557 -1542 -541
rect -1484 -507 -1364 -469
rect -1484 -541 -1468 -507
rect -1380 -541 -1364 -507
rect -1484 -557 -1364 -541
rect -1306 -507 -1186 -469
rect -1306 -541 -1290 -507
rect -1202 -541 -1186 -507
rect -1306 -557 -1186 -541
rect -1128 -507 -1008 -469
rect -1128 -541 -1112 -507
rect -1024 -541 -1008 -507
rect -1128 -557 -1008 -541
rect -950 -507 -830 -469
rect -950 -541 -934 -507
rect -846 -541 -830 -507
rect -950 -557 -830 -541
rect -772 -507 -652 -469
rect -772 -541 -756 -507
rect -668 -541 -652 -507
rect -772 -557 -652 -541
rect -594 -507 -474 -469
rect -594 -541 -578 -507
rect -490 -541 -474 -507
rect -594 -557 -474 -541
rect -416 -507 -296 -469
rect -416 -541 -400 -507
rect -312 -541 -296 -507
rect -416 -557 -296 -541
rect -238 -507 -118 -469
rect -238 -541 -222 -507
rect -134 -541 -118 -507
rect -238 -557 -118 -541
rect -60 -507 60 -469
rect -60 -541 -44 -507
rect 44 -541 60 -507
rect -60 -557 60 -541
rect 118 -507 238 -469
rect 118 -541 134 -507
rect 222 -541 238 -507
rect 118 -557 238 -541
rect 296 -507 416 -469
rect 296 -541 312 -507
rect 400 -541 416 -507
rect 296 -557 416 -541
rect 474 -507 594 -469
rect 474 -541 490 -507
rect 578 -541 594 -507
rect 474 -557 594 -541
rect 652 -507 772 -469
rect 652 -541 668 -507
rect 756 -541 772 -507
rect 652 -557 772 -541
rect 830 -507 950 -469
rect 830 -541 846 -507
rect 934 -541 950 -507
rect 830 -557 950 -541
rect 1008 -507 1128 -469
rect 1008 -541 1024 -507
rect 1112 -541 1128 -507
rect 1008 -557 1128 -541
rect 1186 -507 1306 -469
rect 1186 -541 1202 -507
rect 1290 -541 1306 -507
rect 1186 -557 1306 -541
rect 1364 -507 1484 -469
rect 1364 -541 1380 -507
rect 1468 -541 1484 -507
rect 1364 -557 1484 -541
rect 1542 -507 1662 -469
rect 1542 -541 1558 -507
rect 1646 -541 1662 -507
rect 1542 -557 1662 -541
rect 1720 -507 1840 -469
rect 1720 -541 1736 -507
rect 1824 -541 1840 -507
rect 1720 -557 1840 -541
rect 1898 -507 2018 -469
rect 1898 -541 1914 -507
rect 2002 -541 2018 -507
rect 1898 -557 2018 -541
rect 2076 -507 2196 -469
rect 2076 -541 2092 -507
rect 2180 -541 2196 -507
rect 2076 -557 2196 -541
rect 2254 -507 2374 -469
rect 2254 -541 2270 -507
rect 2358 -541 2374 -507
rect 2254 -557 2374 -541
rect 2432 -507 2552 -469
rect 2432 -541 2448 -507
rect 2536 -541 2552 -507
rect 2432 -557 2552 -541
rect 2610 -507 2730 -469
rect 2610 -541 2626 -507
rect 2714 -541 2730 -507
rect 2610 -557 2730 -541
rect 2788 -507 2908 -469
rect 2788 -541 2804 -507
rect 2892 -541 2908 -507
rect 2788 -557 2908 -541
rect 2966 -507 3086 -469
rect 2966 -541 2982 -507
rect 3070 -541 3086 -507
rect 2966 -557 3086 -541
rect 3144 -507 3264 -469
rect 3144 -541 3160 -507
rect 3248 -541 3264 -507
rect 3144 -557 3264 -541
rect 3322 -507 3442 -469
rect 3322 -541 3338 -507
rect 3426 -541 3442 -507
rect 3322 -557 3442 -541
rect 3500 -507 3620 -469
rect 3500 -541 3516 -507
rect 3604 -541 3620 -507
rect 3500 -557 3620 -541
rect 3678 -507 3798 -469
rect 3678 -541 3694 -507
rect 3782 -541 3798 -507
rect 3678 -557 3798 -541
rect 3856 -507 3976 -469
rect 3856 -541 3872 -507
rect 3960 -541 3976 -507
rect 3856 -557 3976 -541
rect 4034 -507 4154 -469
rect 4034 -541 4050 -507
rect 4138 -541 4154 -507
rect 4034 -557 4154 -541
<< polycont >>
rect -4138 -541 -4050 -507
rect -3960 -541 -3872 -507
rect -3782 -541 -3694 -507
rect -3604 -541 -3516 -507
rect -3426 -541 -3338 -507
rect -3248 -541 -3160 -507
rect -3070 -541 -2982 -507
rect -2892 -541 -2804 -507
rect -2714 -541 -2626 -507
rect -2536 -541 -2448 -507
rect -2358 -541 -2270 -507
rect -2180 -541 -2092 -507
rect -2002 -541 -1914 -507
rect -1824 -541 -1736 -507
rect -1646 -541 -1558 -507
rect -1468 -541 -1380 -507
rect -1290 -541 -1202 -507
rect -1112 -541 -1024 -507
rect -934 -541 -846 -507
rect -756 -541 -668 -507
rect -578 -541 -490 -507
rect -400 -541 -312 -507
rect -222 -541 -134 -507
rect -44 -541 44 -507
rect 134 -541 222 -507
rect 312 -541 400 -507
rect 490 -541 578 -507
rect 668 -541 756 -507
rect 846 -541 934 -507
rect 1024 -541 1112 -507
rect 1202 -541 1290 -507
rect 1380 -541 1468 -507
rect 1558 -541 1646 -507
rect 1736 -541 1824 -507
rect 1914 -541 2002 -507
rect 2092 -541 2180 -507
rect 2270 -541 2358 -507
rect 2448 -541 2536 -507
rect 2626 -541 2714 -507
rect 2804 -541 2892 -507
rect 2982 -541 3070 -507
rect 3160 -541 3248 -507
rect 3338 -541 3426 -507
rect 3516 -541 3604 -507
rect 3694 -541 3782 -507
rect 3872 -541 3960 -507
rect 4050 -541 4138 -507
<< locali >>
rect -4334 645 -4238 679
rect 4238 645 4334 679
rect -4334 583 -4300 645
rect 4300 583 4334 645
rect -4200 519 -4166 535
rect -4200 -473 -4166 -457
rect -4022 519 -3988 535
rect -4022 -473 -3988 -457
rect -3844 519 -3810 535
rect -3844 -473 -3810 -457
rect -3666 519 -3632 535
rect -3666 -473 -3632 -457
rect -3488 519 -3454 535
rect -3488 -473 -3454 -457
rect -3310 519 -3276 535
rect -3310 -473 -3276 -457
rect -3132 519 -3098 535
rect -3132 -473 -3098 -457
rect -2954 519 -2920 535
rect -2954 -473 -2920 -457
rect -2776 519 -2742 535
rect -2776 -473 -2742 -457
rect -2598 519 -2564 535
rect -2598 -473 -2564 -457
rect -2420 519 -2386 535
rect -2420 -473 -2386 -457
rect -2242 519 -2208 535
rect -2242 -473 -2208 -457
rect -2064 519 -2030 535
rect -2064 -473 -2030 -457
rect -1886 519 -1852 535
rect -1886 -473 -1852 -457
rect -1708 519 -1674 535
rect -1708 -473 -1674 -457
rect -1530 519 -1496 535
rect -1530 -473 -1496 -457
rect -1352 519 -1318 535
rect -1352 -473 -1318 -457
rect -1174 519 -1140 535
rect -1174 -473 -1140 -457
rect -996 519 -962 535
rect -996 -473 -962 -457
rect -818 519 -784 535
rect -818 -473 -784 -457
rect -640 519 -606 535
rect -640 -473 -606 -457
rect -462 519 -428 535
rect -462 -473 -428 -457
rect -284 519 -250 535
rect -284 -473 -250 -457
rect -106 519 -72 535
rect -106 -473 -72 -457
rect 72 519 106 535
rect 72 -473 106 -457
rect 250 519 284 535
rect 250 -473 284 -457
rect 428 519 462 535
rect 428 -473 462 -457
rect 606 519 640 535
rect 606 -473 640 -457
rect 784 519 818 535
rect 784 -473 818 -457
rect 962 519 996 535
rect 962 -473 996 -457
rect 1140 519 1174 535
rect 1140 -473 1174 -457
rect 1318 519 1352 535
rect 1318 -473 1352 -457
rect 1496 519 1530 535
rect 1496 -473 1530 -457
rect 1674 519 1708 535
rect 1674 -473 1708 -457
rect 1852 519 1886 535
rect 1852 -473 1886 -457
rect 2030 519 2064 535
rect 2030 -473 2064 -457
rect 2208 519 2242 535
rect 2208 -473 2242 -457
rect 2386 519 2420 535
rect 2386 -473 2420 -457
rect 2564 519 2598 535
rect 2564 -473 2598 -457
rect 2742 519 2776 535
rect 2742 -473 2776 -457
rect 2920 519 2954 535
rect 2920 -473 2954 -457
rect 3098 519 3132 535
rect 3098 -473 3132 -457
rect 3276 519 3310 535
rect 3276 -473 3310 -457
rect 3454 519 3488 535
rect 3454 -473 3488 -457
rect 3632 519 3666 535
rect 3632 -473 3666 -457
rect 3810 519 3844 535
rect 3810 -473 3844 -457
rect 3988 519 4022 535
rect 3988 -473 4022 -457
rect 4166 519 4200 535
rect 4166 -473 4200 -457
rect -4154 -541 -4138 -507
rect -4050 -541 -4034 -507
rect -3976 -541 -3960 -507
rect -3872 -541 -3856 -507
rect -3798 -541 -3782 -507
rect -3694 -541 -3678 -507
rect -3620 -541 -3604 -507
rect -3516 -541 -3500 -507
rect -3442 -541 -3426 -507
rect -3338 -541 -3322 -507
rect -3264 -541 -3248 -507
rect -3160 -541 -3144 -507
rect -3086 -541 -3070 -507
rect -2982 -541 -2966 -507
rect -2908 -541 -2892 -507
rect -2804 -541 -2788 -507
rect -2730 -541 -2714 -507
rect -2626 -541 -2610 -507
rect -2552 -541 -2536 -507
rect -2448 -541 -2432 -507
rect -2374 -541 -2358 -507
rect -2270 -541 -2254 -507
rect -2196 -541 -2180 -507
rect -2092 -541 -2076 -507
rect -2018 -541 -2002 -507
rect -1914 -541 -1898 -507
rect -1840 -541 -1824 -507
rect -1736 -541 -1720 -507
rect -1662 -541 -1646 -507
rect -1558 -541 -1542 -507
rect -1484 -541 -1468 -507
rect -1380 -541 -1364 -507
rect -1306 -541 -1290 -507
rect -1202 -541 -1186 -507
rect -1128 -541 -1112 -507
rect -1024 -541 -1008 -507
rect -950 -541 -934 -507
rect -846 -541 -830 -507
rect -772 -541 -756 -507
rect -668 -541 -652 -507
rect -594 -541 -578 -507
rect -490 -541 -474 -507
rect -416 -541 -400 -507
rect -312 -541 -296 -507
rect -238 -541 -222 -507
rect -134 -541 -118 -507
rect -60 -541 -44 -507
rect 44 -541 60 -507
rect 118 -541 134 -507
rect 222 -541 238 -507
rect 296 -541 312 -507
rect 400 -541 416 -507
rect 474 -541 490 -507
rect 578 -541 594 -507
rect 652 -541 668 -507
rect 756 -541 772 -507
rect 830 -541 846 -507
rect 934 -541 950 -507
rect 1008 -541 1024 -507
rect 1112 -541 1128 -507
rect 1186 -541 1202 -507
rect 1290 -541 1306 -507
rect 1364 -541 1380 -507
rect 1468 -541 1484 -507
rect 1542 -541 1558 -507
rect 1646 -541 1662 -507
rect 1720 -541 1736 -507
rect 1824 -541 1840 -507
rect 1898 -541 1914 -507
rect 2002 -541 2018 -507
rect 2076 -541 2092 -507
rect 2180 -541 2196 -507
rect 2254 -541 2270 -507
rect 2358 -541 2374 -507
rect 2432 -541 2448 -507
rect 2536 -541 2552 -507
rect 2610 -541 2626 -507
rect 2714 -541 2730 -507
rect 2788 -541 2804 -507
rect 2892 -541 2908 -507
rect 2966 -541 2982 -507
rect 3070 -541 3086 -507
rect 3144 -541 3160 -507
rect 3248 -541 3264 -507
rect 3322 -541 3338 -507
rect 3426 -541 3442 -507
rect 3500 -541 3516 -507
rect 3604 -541 3620 -507
rect 3678 -541 3694 -507
rect 3782 -541 3798 -507
rect 3856 -541 3872 -507
rect 3960 -541 3976 -507
rect 4034 -541 4050 -507
rect 4138 -541 4154 -507
rect -4334 -645 -4300 -583
rect 4300 -645 4334 -583
rect -4334 -679 -4238 -645
rect 4238 -679 4334 -645
<< viali >>
rect -4200 -457 -4166 519
rect -4022 -457 -3988 519
rect -3844 -457 -3810 519
rect -3666 -457 -3632 519
rect -3488 -457 -3454 519
rect -3310 -457 -3276 519
rect -3132 -457 -3098 519
rect -2954 -457 -2920 519
rect -2776 -457 -2742 519
rect -2598 -457 -2564 519
rect -2420 -457 -2386 519
rect -2242 -457 -2208 519
rect -2064 -457 -2030 519
rect -1886 -457 -1852 519
rect -1708 -457 -1674 519
rect -1530 -457 -1496 519
rect -1352 -457 -1318 519
rect -1174 -457 -1140 519
rect -996 -457 -962 519
rect -818 -457 -784 519
rect -640 -457 -606 519
rect -462 -457 -428 519
rect -284 -457 -250 519
rect -106 -457 -72 519
rect 72 -457 106 519
rect 250 -457 284 519
rect 428 -457 462 519
rect 606 -457 640 519
rect 784 -457 818 519
rect 962 -457 996 519
rect 1140 -457 1174 519
rect 1318 -457 1352 519
rect 1496 -457 1530 519
rect 1674 -457 1708 519
rect 1852 -457 1886 519
rect 2030 -457 2064 519
rect 2208 -457 2242 519
rect 2386 -457 2420 519
rect 2564 -457 2598 519
rect 2742 -457 2776 519
rect 2920 -457 2954 519
rect 3098 -457 3132 519
rect 3276 -457 3310 519
rect 3454 -457 3488 519
rect 3632 -457 3666 519
rect 3810 -457 3844 519
rect 3988 -457 4022 519
rect 4166 -457 4200 519
rect -4138 -541 -4050 -507
rect -3960 -541 -3872 -507
rect -3782 -541 -3694 -507
rect -3604 -541 -3516 -507
rect -3426 -541 -3338 -507
rect -3248 -541 -3160 -507
rect -3070 -541 -2982 -507
rect -2892 -541 -2804 -507
rect -2714 -541 -2626 -507
rect -2536 -541 -2448 -507
rect -2358 -541 -2270 -507
rect -2180 -541 -2092 -507
rect -2002 -541 -1914 -507
rect -1824 -541 -1736 -507
rect -1646 -541 -1558 -507
rect -1468 -541 -1380 -507
rect -1290 -541 -1202 -507
rect -1112 -541 -1024 -507
rect -934 -541 -846 -507
rect -756 -541 -668 -507
rect -578 -541 -490 -507
rect -400 -541 -312 -507
rect -222 -541 -134 -507
rect -44 -541 44 -507
rect 134 -541 222 -507
rect 312 -541 400 -507
rect 490 -541 578 -507
rect 668 -541 756 -507
rect 846 -541 934 -507
rect 1024 -541 1112 -507
rect 1202 -541 1290 -507
rect 1380 -541 1468 -507
rect 1558 -541 1646 -507
rect 1736 -541 1824 -507
rect 1914 -541 2002 -507
rect 2092 -541 2180 -507
rect 2270 -541 2358 -507
rect 2448 -541 2536 -507
rect 2626 -541 2714 -507
rect 2804 -541 2892 -507
rect 2982 -541 3070 -507
rect 3160 -541 3248 -507
rect 3338 -541 3426 -507
rect 3516 -541 3604 -507
rect 3694 -541 3782 -507
rect 3872 -541 3960 -507
rect 4050 -541 4138 -507
<< metal1 >>
rect -4206 519 -4160 531
rect -4206 -457 -4200 519
rect -4166 -457 -4160 519
rect -4206 -469 -4160 -457
rect -4028 519 -3982 531
rect -4028 -457 -4022 519
rect -3988 -457 -3982 519
rect -4028 -469 -3982 -457
rect -3850 519 -3804 531
rect -3850 -457 -3844 519
rect -3810 -457 -3804 519
rect -3850 -469 -3804 -457
rect -3672 519 -3626 531
rect -3672 -457 -3666 519
rect -3632 -457 -3626 519
rect -3672 -469 -3626 -457
rect -3494 519 -3448 531
rect -3494 -457 -3488 519
rect -3454 -457 -3448 519
rect -3494 -469 -3448 -457
rect -3316 519 -3270 531
rect -3316 -457 -3310 519
rect -3276 -457 -3270 519
rect -3316 -469 -3270 -457
rect -3138 519 -3092 531
rect -3138 -457 -3132 519
rect -3098 -457 -3092 519
rect -3138 -469 -3092 -457
rect -2960 519 -2914 531
rect -2960 -457 -2954 519
rect -2920 -457 -2914 519
rect -2960 -469 -2914 -457
rect -2782 519 -2736 531
rect -2782 -457 -2776 519
rect -2742 -457 -2736 519
rect -2782 -469 -2736 -457
rect -2604 519 -2558 531
rect -2604 -457 -2598 519
rect -2564 -457 -2558 519
rect -2604 -469 -2558 -457
rect -2426 519 -2380 531
rect -2426 -457 -2420 519
rect -2386 -457 -2380 519
rect -2426 -469 -2380 -457
rect -2248 519 -2202 531
rect -2248 -457 -2242 519
rect -2208 -457 -2202 519
rect -2248 -469 -2202 -457
rect -2070 519 -2024 531
rect -2070 -457 -2064 519
rect -2030 -457 -2024 519
rect -2070 -469 -2024 -457
rect -1892 519 -1846 531
rect -1892 -457 -1886 519
rect -1852 -457 -1846 519
rect -1892 -469 -1846 -457
rect -1714 519 -1668 531
rect -1714 -457 -1708 519
rect -1674 -457 -1668 519
rect -1714 -469 -1668 -457
rect -1536 519 -1490 531
rect -1536 -457 -1530 519
rect -1496 -457 -1490 519
rect -1536 -469 -1490 -457
rect -1358 519 -1312 531
rect -1358 -457 -1352 519
rect -1318 -457 -1312 519
rect -1358 -469 -1312 -457
rect -1180 519 -1134 531
rect -1180 -457 -1174 519
rect -1140 -457 -1134 519
rect -1180 -469 -1134 -457
rect -1002 519 -956 531
rect -1002 -457 -996 519
rect -962 -457 -956 519
rect -1002 -469 -956 -457
rect -824 519 -778 531
rect -824 -457 -818 519
rect -784 -457 -778 519
rect -824 -469 -778 -457
rect -646 519 -600 531
rect -646 -457 -640 519
rect -606 -457 -600 519
rect -646 -469 -600 -457
rect -468 519 -422 531
rect -468 -457 -462 519
rect -428 -457 -422 519
rect -468 -469 -422 -457
rect -290 519 -244 531
rect -290 -457 -284 519
rect -250 -457 -244 519
rect -290 -469 -244 -457
rect -112 519 -66 531
rect -112 -457 -106 519
rect -72 -457 -66 519
rect -112 -469 -66 -457
rect 66 519 112 531
rect 66 -457 72 519
rect 106 -457 112 519
rect 66 -469 112 -457
rect 244 519 290 531
rect 244 -457 250 519
rect 284 -457 290 519
rect 244 -469 290 -457
rect 422 519 468 531
rect 422 -457 428 519
rect 462 -457 468 519
rect 422 -469 468 -457
rect 600 519 646 531
rect 600 -457 606 519
rect 640 -457 646 519
rect 600 -469 646 -457
rect 778 519 824 531
rect 778 -457 784 519
rect 818 -457 824 519
rect 778 -469 824 -457
rect 956 519 1002 531
rect 956 -457 962 519
rect 996 -457 1002 519
rect 956 -469 1002 -457
rect 1134 519 1180 531
rect 1134 -457 1140 519
rect 1174 -457 1180 519
rect 1134 -469 1180 -457
rect 1312 519 1358 531
rect 1312 -457 1318 519
rect 1352 -457 1358 519
rect 1312 -469 1358 -457
rect 1490 519 1536 531
rect 1490 -457 1496 519
rect 1530 -457 1536 519
rect 1490 -469 1536 -457
rect 1668 519 1714 531
rect 1668 -457 1674 519
rect 1708 -457 1714 519
rect 1668 -469 1714 -457
rect 1846 519 1892 531
rect 1846 -457 1852 519
rect 1886 -457 1892 519
rect 1846 -469 1892 -457
rect 2024 519 2070 531
rect 2024 -457 2030 519
rect 2064 -457 2070 519
rect 2024 -469 2070 -457
rect 2202 519 2248 531
rect 2202 -457 2208 519
rect 2242 -457 2248 519
rect 2202 -469 2248 -457
rect 2380 519 2426 531
rect 2380 -457 2386 519
rect 2420 -457 2426 519
rect 2380 -469 2426 -457
rect 2558 519 2604 531
rect 2558 -457 2564 519
rect 2598 -457 2604 519
rect 2558 -469 2604 -457
rect 2736 519 2782 531
rect 2736 -457 2742 519
rect 2776 -457 2782 519
rect 2736 -469 2782 -457
rect 2914 519 2960 531
rect 2914 -457 2920 519
rect 2954 -457 2960 519
rect 2914 -469 2960 -457
rect 3092 519 3138 531
rect 3092 -457 3098 519
rect 3132 -457 3138 519
rect 3092 -469 3138 -457
rect 3270 519 3316 531
rect 3270 -457 3276 519
rect 3310 -457 3316 519
rect 3270 -469 3316 -457
rect 3448 519 3494 531
rect 3448 -457 3454 519
rect 3488 -457 3494 519
rect 3448 -469 3494 -457
rect 3626 519 3672 531
rect 3626 -457 3632 519
rect 3666 -457 3672 519
rect 3626 -469 3672 -457
rect 3804 519 3850 531
rect 3804 -457 3810 519
rect 3844 -457 3850 519
rect 3804 -469 3850 -457
rect 3982 519 4028 531
rect 3982 -457 3988 519
rect 4022 -457 4028 519
rect 3982 -469 4028 -457
rect 4160 519 4206 531
rect 4160 -457 4166 519
rect 4200 -457 4206 519
rect 4160 -469 4206 -457
rect -4150 -507 -4038 -501
rect -4150 -541 -4138 -507
rect -4050 -541 -4038 -507
rect -4150 -547 -4038 -541
rect -3972 -507 -3860 -501
rect -3972 -541 -3960 -507
rect -3872 -541 -3860 -507
rect -3972 -547 -3860 -541
rect -3794 -507 -3682 -501
rect -3794 -541 -3782 -507
rect -3694 -541 -3682 -507
rect -3794 -547 -3682 -541
rect -3616 -507 -3504 -501
rect -3616 -541 -3604 -507
rect -3516 -541 -3504 -507
rect -3616 -547 -3504 -541
rect -3438 -507 -3326 -501
rect -3438 -541 -3426 -507
rect -3338 -541 -3326 -507
rect -3438 -547 -3326 -541
rect -3260 -507 -3148 -501
rect -3260 -541 -3248 -507
rect -3160 -541 -3148 -507
rect -3260 -547 -3148 -541
rect -3082 -507 -2970 -501
rect -3082 -541 -3070 -507
rect -2982 -541 -2970 -507
rect -3082 -547 -2970 -541
rect -2904 -507 -2792 -501
rect -2904 -541 -2892 -507
rect -2804 -541 -2792 -507
rect -2904 -547 -2792 -541
rect -2726 -507 -2614 -501
rect -2726 -541 -2714 -507
rect -2626 -541 -2614 -507
rect -2726 -547 -2614 -541
rect -2548 -507 -2436 -501
rect -2548 -541 -2536 -507
rect -2448 -541 -2436 -507
rect -2548 -547 -2436 -541
rect -2370 -507 -2258 -501
rect -2370 -541 -2358 -507
rect -2270 -541 -2258 -507
rect -2370 -547 -2258 -541
rect -2192 -507 -2080 -501
rect -2192 -541 -2180 -507
rect -2092 -541 -2080 -507
rect -2192 -547 -2080 -541
rect -2014 -507 -1902 -501
rect -2014 -541 -2002 -507
rect -1914 -541 -1902 -507
rect -2014 -547 -1902 -541
rect -1836 -507 -1724 -501
rect -1836 -541 -1824 -507
rect -1736 -541 -1724 -507
rect -1836 -547 -1724 -541
rect -1658 -507 -1546 -501
rect -1658 -541 -1646 -507
rect -1558 -541 -1546 -507
rect -1658 -547 -1546 -541
rect -1480 -507 -1368 -501
rect -1480 -541 -1468 -507
rect -1380 -541 -1368 -507
rect -1480 -547 -1368 -541
rect -1302 -507 -1190 -501
rect -1302 -541 -1290 -507
rect -1202 -541 -1190 -507
rect -1302 -547 -1190 -541
rect -1124 -507 -1012 -501
rect -1124 -541 -1112 -507
rect -1024 -541 -1012 -507
rect -1124 -547 -1012 -541
rect -946 -507 -834 -501
rect -946 -541 -934 -507
rect -846 -541 -834 -507
rect -946 -547 -834 -541
rect -768 -507 -656 -501
rect -768 -541 -756 -507
rect -668 -541 -656 -507
rect -768 -547 -656 -541
rect -590 -507 -478 -501
rect -590 -541 -578 -507
rect -490 -541 -478 -507
rect -590 -547 -478 -541
rect -412 -507 -300 -501
rect -412 -541 -400 -507
rect -312 -541 -300 -507
rect -412 -547 -300 -541
rect -234 -507 -122 -501
rect -234 -541 -222 -507
rect -134 -541 -122 -507
rect -234 -547 -122 -541
rect -56 -507 56 -501
rect -56 -541 -44 -507
rect 44 -541 56 -507
rect -56 -547 56 -541
rect 122 -507 234 -501
rect 122 -541 134 -507
rect 222 -541 234 -507
rect 122 -547 234 -541
rect 300 -507 412 -501
rect 300 -541 312 -507
rect 400 -541 412 -507
rect 300 -547 412 -541
rect 478 -507 590 -501
rect 478 -541 490 -507
rect 578 -541 590 -507
rect 478 -547 590 -541
rect 656 -507 768 -501
rect 656 -541 668 -507
rect 756 -541 768 -507
rect 656 -547 768 -541
rect 834 -507 946 -501
rect 834 -541 846 -507
rect 934 -541 946 -507
rect 834 -547 946 -541
rect 1012 -507 1124 -501
rect 1012 -541 1024 -507
rect 1112 -541 1124 -507
rect 1012 -547 1124 -541
rect 1190 -507 1302 -501
rect 1190 -541 1202 -507
rect 1290 -541 1302 -507
rect 1190 -547 1302 -541
rect 1368 -507 1480 -501
rect 1368 -541 1380 -507
rect 1468 -541 1480 -507
rect 1368 -547 1480 -541
rect 1546 -507 1658 -501
rect 1546 -541 1558 -507
rect 1646 -541 1658 -507
rect 1546 -547 1658 -541
rect 1724 -507 1836 -501
rect 1724 -541 1736 -507
rect 1824 -541 1836 -507
rect 1724 -547 1836 -541
rect 1902 -507 2014 -501
rect 1902 -541 1914 -507
rect 2002 -541 2014 -507
rect 1902 -547 2014 -541
rect 2080 -507 2192 -501
rect 2080 -541 2092 -507
rect 2180 -541 2192 -507
rect 2080 -547 2192 -541
rect 2258 -507 2370 -501
rect 2258 -541 2270 -507
rect 2358 -541 2370 -507
rect 2258 -547 2370 -541
rect 2436 -507 2548 -501
rect 2436 -541 2448 -507
rect 2536 -541 2548 -507
rect 2436 -547 2548 -541
rect 2614 -507 2726 -501
rect 2614 -541 2626 -507
rect 2714 -541 2726 -507
rect 2614 -547 2726 -541
rect 2792 -507 2904 -501
rect 2792 -541 2804 -507
rect 2892 -541 2904 -507
rect 2792 -547 2904 -541
rect 2970 -507 3082 -501
rect 2970 -541 2982 -507
rect 3070 -541 3082 -507
rect 2970 -547 3082 -541
rect 3148 -507 3260 -501
rect 3148 -541 3160 -507
rect 3248 -541 3260 -507
rect 3148 -547 3260 -541
rect 3326 -507 3438 -501
rect 3326 -541 3338 -507
rect 3426 -541 3438 -507
rect 3326 -547 3438 -541
rect 3504 -507 3616 -501
rect 3504 -541 3516 -507
rect 3604 -541 3616 -507
rect 3504 -547 3616 -541
rect 3682 -507 3794 -501
rect 3682 -541 3694 -507
rect 3782 -541 3794 -507
rect 3682 -547 3794 -541
rect 3860 -507 3972 -501
rect 3860 -541 3872 -507
rect 3960 -541 3972 -507
rect 3860 -547 3972 -541
rect 4038 -507 4150 -501
rect 4038 -541 4050 -507
rect 4138 -541 4150 -507
rect 4038 -547 4150 -541
<< properties >>
string FIXED_BBOX -4317 -662 4317 662
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.6 m 1 nf 47 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
