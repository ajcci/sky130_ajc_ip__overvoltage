magic
tech sky130A
magscale 1 2
timestamp 1712627826
<< nwell >>
rect 13226 11244 13282 11290
rect 13236 10162 13282 10205
rect 10168 9524 13488 9906
<< pwell >>
rect 1224 8514 1270 8546
rect 7220 8468 7276 8514
<< locali >>
rect 1078 10697 1142 10712
rect 1078 10599 1093 10697
rect 1127 10599 1142 10697
rect 1078 10584 1142 10599
rect 13360 10697 13424 10712
rect 13360 10599 13375 10697
rect 13409 10599 13424 10697
rect 13360 10584 13424 10599
rect 1078 9197 1142 9212
rect 1078 9099 1093 9197
rect 1127 9099 1142 9197
rect 1078 9084 1142 9099
rect 7355 9197 7419 9212
rect 7355 9099 7370 9197
rect 7404 9099 7419 9197
rect 7355 9084 7419 9099
rect 10231 8662 10295 8677
rect 10231 8564 10246 8662
rect 10280 8564 10295 8662
rect 10231 8549 10295 8564
rect 12099 8662 12163 8677
rect 12099 8564 12114 8662
rect 12148 8564 12163 8662
rect 12099 8549 12163 8564
rect 14659 8662 14723 8677
rect 14659 8564 14674 8662
rect 14708 8564 14723 8662
rect 14659 8549 14723 8564
rect 115 8075 243 8090
rect 7643 8060 7707 8075
rect 115 8026 243 8041
rect 7643 7962 7658 8060
rect 7692 7962 7707 8060
rect 15112 8042 15312 8146
rect 7643 7947 7707 7962
rect 15112 7621 15296 7725
rect 8857 6839 8921 6854
rect 8857 6741 8872 6839
rect 8906 6741 8921 6839
rect 8857 6726 8921 6741
rect 12151 6839 12215 6854
rect 12151 6741 12166 6839
rect 12200 6741 12215 6839
rect 12151 6726 12215 6741
rect 12319 6839 12383 6854
rect 12319 6741 12334 6839
rect 12368 6741 12383 6839
rect 12319 6726 12383 6741
rect 14418 6839 14482 6854
rect 14418 6741 14433 6839
rect 14467 6741 14482 6839
rect 14418 6726 14482 6741
rect 15112 6373 15312 6477
rect 8483 5526 8498 5654
rect 8483 4370 8498 4498
rect 8483 3214 8498 3342
rect 8483 2058 8498 2186
rect 8483 902 8498 1030
rect 7643 96 7673 111
rect 7643 -2 7658 96
rect 8532 5526 8547 5654
rect 15383 5526 15398 5654
rect 8532 4370 8547 4498
rect 15383 4370 15398 4498
rect 8532 3214 8547 3342
rect 15383 3214 15398 3342
rect 8532 2058 8547 2186
rect 15383 2058 15398 2186
rect 8532 902 8547 1030
rect 15383 902 15398 1030
rect 15432 5526 15447 5654
rect 15432 4370 15447 4498
rect 15432 3214 15447 3342
rect 15432 2058 15447 2186
rect 15432 902 15447 1030
rect 7692 -2 7707 79
rect 7643 -17 7707 -2
<< viali >>
rect 1192 11388 13314 11422
rect 1093 10599 1127 10697
rect 13375 10599 13409 10697
rect 1192 9984 13314 10018
rect 1192 9722 7308 9756
rect 10342 9412 15654 9446
rect 1093 9099 1127 9197
rect 7370 9099 7404 9197
rect 10246 8564 10280 8662
rect 12114 8564 12148 8662
rect 14674 8564 14708 8662
rect 1192 8336 7308 8370
rect 79 8041 7611 8075
rect -17 79 17 7979
rect 7658 7962 7692 8060
rect 10342 8008 15654 8042
rect 7673 148 7707 7911
rect 8872 6741 8906 6839
rect 12166 6741 12200 6839
rect 12334 6741 12368 6839
rect 14433 6741 14467 6839
rect 8594 5931 15336 5965
rect 79 -17 7611 17
rect 7658 -2 7692 96
rect 8498 79 8532 5869
rect 15398 79 15432 5869
rect 8594 -17 15336 17
<< metal1 >>
rect 1084 11422 13422 11434
rect 1084 11388 1192 11422
rect 13314 11388 13422 11422
rect 1084 11376 13422 11388
rect 1084 10722 1142 11376
rect 3640 11307 3788 11318
rect 1224 11244 1280 11290
rect 2930 11244 2996 11290
rect 3640 11255 3651 11307
rect 3777 11255 3788 11307
rect 3640 11244 3788 11255
rect 4712 11307 4860 11318
rect 4712 11255 4723 11307
rect 4849 11255 4860 11307
rect 7172 11290 7220 11376
rect 4712 11244 4860 11255
rect 5504 11244 5570 11290
rect 8078 11244 8144 11290
rect 8936 11244 9002 11290
rect 9794 11244 9860 11290
rect 11510 11244 11576 11290
rect 13226 11244 13282 11290
rect 1224 11203 1270 11244
rect 4600 11203 4646 11244
rect 5514 11203 5560 11244
rect 7172 11203 7220 11244
rect 11520 11203 11566 11244
rect 13236 11203 13282 11244
rect 4600 11157 4656 11203
rect 7172 11155 7230 11203
rect 8074 11192 8148 11203
rect 8074 11066 8085 11192
rect 8137 11066 8148 11192
rect 8074 11055 8148 11066
rect 9790 11192 9864 11203
rect 9790 11066 9801 11192
rect 9853 11066 9864 11192
rect 9790 11055 9864 11066
rect 13364 10722 13422 11376
rect 1073 10711 1147 10722
rect 1073 10585 1084 10711
rect 1136 10585 1147 10711
rect 1073 10574 1147 10585
rect 1209 10711 1283 10722
rect 1209 10585 1220 10711
rect 1272 10585 1283 10711
rect 1209 10574 1283 10585
rect 2067 10711 2141 10722
rect 2067 10585 2078 10711
rect 2130 10585 2141 10711
rect 2067 10574 2141 10585
rect 3783 10711 3857 10722
rect 3783 10585 3794 10711
rect 3846 10585 3857 10711
rect 3783 10574 3857 10585
rect 4641 10711 4715 10722
rect 4641 10585 4652 10711
rect 4704 10585 4715 10711
rect 4641 10574 4715 10585
rect 6357 10711 6431 10722
rect 6357 10585 6368 10711
rect 6420 10585 6431 10711
rect 6357 10574 6431 10585
rect 7216 10711 7290 10722
rect 7216 10585 7227 10711
rect 7279 10585 7290 10711
rect 7216 10574 7290 10585
rect 8932 10711 9006 10722
rect 8932 10585 8943 10711
rect 8995 10585 9006 10711
rect 8932 10574 9006 10585
rect 10648 10711 10722 10722
rect 10648 10585 10659 10711
rect 10711 10585 10722 10711
rect 10648 10574 10722 10585
rect 12364 10711 12438 10722
rect 12364 10585 12375 10711
rect 12427 10585 12438 10711
rect 12364 10574 12438 10585
rect 13222 10711 13296 10722
rect 13222 10585 13233 10711
rect 13285 10585 13296 10711
rect 13222 10574 13296 10585
rect 13355 10711 13429 10722
rect 13355 10585 13366 10711
rect 13418 10585 13429 10711
rect 13355 10574 13429 10585
rect 1084 10030 1142 10574
rect 2931 10325 2995 10331
rect 2931 10209 2937 10325
rect 2989 10209 2995 10325
rect 5505 10325 5569 10331
rect 2931 10203 2995 10209
rect 4600 10203 4656 10249
rect 5505 10209 5511 10325
rect 5563 10209 5569 10325
rect 1224 10162 1270 10203
rect 4600 10162 4646 10203
rect 5505 10162 5569 10209
rect 7172 10203 7230 10251
rect 1224 10116 1280 10162
rect 2930 10116 2996 10162
rect 3640 10151 3788 10162
rect 3640 10099 3651 10151
rect 3777 10099 3788 10151
rect 3640 10088 3788 10099
rect 4712 10151 4860 10162
rect 4712 10099 4723 10151
rect 4849 10099 4860 10151
rect 5504 10116 5570 10162
rect 4712 10088 4860 10099
rect 7172 10030 7220 10203
rect 11520 10189 11566 10203
rect 11427 10183 11566 10189
rect 10255 10172 10383 10178
rect 8078 10116 8144 10162
rect 8936 10116 9002 10162
rect 9794 10116 9860 10162
rect 10255 10120 10261 10172
rect 10377 10120 10383 10172
rect 11427 10131 11433 10183
rect 11549 10162 11566 10183
rect 13236 10162 13282 10205
rect 11549 10131 11576 10162
rect 11427 10125 11576 10131
rect 10255 10114 10383 10120
rect 11510 10116 11576 10125
rect 13226 10116 13282 10162
rect 13364 10030 13422 10574
rect 1084 10018 13422 10030
rect 1084 9984 1192 10018
rect 13314 9984 13422 10018
rect 1084 9972 13422 9984
rect 1084 9756 7416 9768
rect 1084 9722 1192 9756
rect 7308 9722 7416 9756
rect 1084 9710 7416 9722
rect 1084 9222 1142 9710
rect 3640 9647 3788 9658
rect 1224 9578 1280 9624
rect 2930 9578 2996 9624
rect 3640 9595 3651 9647
rect 3777 9595 3788 9647
rect 3640 9584 3788 9595
rect 4712 9647 4860 9658
rect 4712 9595 4723 9647
rect 4849 9595 4860 9647
rect 4712 9584 4860 9595
rect 5504 9584 5570 9624
rect 7220 9578 7276 9624
rect 1224 9546 1270 9578
rect 2931 9546 2995 9578
rect 7230 9546 7276 9578
rect 2931 9430 2937 9546
rect 2989 9430 2995 9546
rect 2931 9424 2995 9430
rect 5505 9430 5511 9546
rect 5563 9430 5569 9546
rect 5505 9424 5569 9430
rect 7358 9222 7416 9710
rect 10234 9446 15762 9458
rect 10234 9412 10342 9446
rect 15654 9412 15762 9446
rect 10234 9400 15762 9412
rect 1073 9211 1147 9222
rect 1073 9085 1084 9211
rect 1136 9085 1147 9211
rect 1073 9074 1147 9085
rect 1209 9211 1283 9222
rect 1209 9085 1220 9211
rect 1272 9085 1283 9211
rect 7216 9211 7290 9222
rect 1209 9074 1283 9085
rect 4216 9137 4290 9148
rect 4216 9085 4227 9137
rect 4279 9085 4290 9137
rect 1084 8382 1142 9074
rect 2068 8760 2142 8771
rect 2068 8634 2079 8760
rect 2131 8634 2142 8760
rect 2068 8623 2142 8634
rect 3784 8760 3858 8771
rect 3784 8634 3795 8760
rect 3847 8634 3858 8760
rect 3784 8623 3858 8634
rect 1224 8514 1270 8546
rect 2940 8514 2986 8557
rect 4216 8514 4290 9085
rect 7216 9085 7227 9211
rect 7279 9085 7290 9211
rect 7216 9074 7290 9085
rect 7350 9211 7424 9222
rect 7350 9085 7361 9211
rect 7413 9085 7424 9211
rect 7350 9074 7424 9085
rect 4642 8760 4716 8771
rect 4642 8634 4653 8760
rect 4705 8634 4716 8760
rect 4642 8623 4716 8634
rect 6358 8760 6432 8771
rect 6358 8634 6369 8760
rect 6421 8634 6432 8760
rect 6358 8623 6432 8634
rect 7230 8514 7276 8546
rect 1224 8468 1280 8514
rect 2930 8468 2996 8514
rect 3640 8497 3788 8508
rect 3640 8445 3651 8497
rect 3777 8445 3788 8497
rect 3640 8434 3788 8445
rect 4712 8497 4860 8508
rect 4712 8445 4723 8497
rect 4849 8445 4860 8497
rect 5504 8468 5570 8514
rect 7220 8468 7276 8514
rect 4712 8434 4860 8445
rect 7358 8382 7416 9074
rect 10234 8687 10292 9400
rect 10453 9327 10527 9338
rect 10453 9275 10464 9327
rect 10516 9275 10527 9327
rect 10453 9264 10527 9275
rect 10612 9322 10676 9328
rect 10612 9270 10618 9322
rect 10670 9270 10676 9322
rect 11166 9317 11230 9323
rect 10612 9264 10676 9270
rect 10819 9309 10883 9315
rect 10819 9257 10825 9309
rect 10877 9257 10883 9309
rect 11166 9265 11172 9317
rect 11224 9265 11230 9317
rect 11166 9259 11230 9265
rect 11522 9317 11586 9323
rect 11522 9265 11528 9317
rect 11580 9265 11586 9317
rect 11522 9259 11586 9265
rect 11871 9318 11945 9329
rect 11871 9266 11882 9318
rect 11934 9266 11945 9318
rect 10819 9251 10883 9257
rect 11871 9255 11945 9266
rect 12320 9322 12448 9328
rect 12320 9270 12326 9322
rect 12442 9270 12448 9322
rect 12320 9264 12448 9270
rect 13150 9268 13216 9314
rect 13605 9179 13679 9190
rect 10932 9140 11006 9151
rect 10932 9014 10943 9140
rect 10995 9014 11006 9140
rect 13605 9053 13616 9179
rect 13668 9053 13679 9179
rect 13605 9042 13679 9053
rect 10932 9003 11006 9014
rect 12684 9010 12758 9021
rect 11037 8918 11111 8929
rect 11037 8792 11048 8918
rect 11100 8792 11111 8918
rect 12684 8884 12695 9010
rect 12747 8884 12758 9010
rect 12684 8873 12758 8884
rect 14523 8894 14597 8905
rect 11037 8781 11111 8792
rect 11132 8727 11264 8783
rect 14523 8768 14534 8894
rect 14586 8768 14597 8894
rect 14523 8757 14597 8768
rect 10716 8707 10790 8718
rect 10226 8676 10300 8687
rect 10226 8550 10237 8676
rect 10289 8550 10300 8676
rect 10716 8655 10727 8707
rect 10779 8655 10790 8707
rect 15704 8687 15762 9400
rect 10716 8644 10790 8655
rect 12094 8676 12168 8687
rect 10226 8539 10300 8550
rect 12094 8550 12105 8676
rect 12157 8550 12168 8676
rect 12094 8539 12168 8550
rect 12230 8676 12304 8687
rect 12230 8550 12241 8676
rect 12293 8550 12304 8676
rect 12230 8539 12304 8550
rect 13146 8676 13220 8687
rect 13146 8550 13157 8676
rect 13209 8550 13220 8676
rect 13146 8539 13220 8550
rect 14062 8676 14136 8687
rect 14062 8550 14073 8676
rect 14125 8550 14136 8676
rect 14062 8539 14136 8550
rect 14654 8676 14728 8687
rect 14654 8550 14665 8676
rect 14717 8550 14728 8676
rect 14654 8539 14728 8550
rect 14788 8676 14862 8687
rect 14788 8550 14799 8676
rect 14851 8550 14862 8676
rect 14788 8539 14862 8550
rect 15562 8676 15636 8687
rect 15562 8550 15573 8676
rect 15625 8550 15636 8676
rect 15562 8539 15636 8550
rect 15694 8676 15768 8687
rect 15694 8550 15705 8676
rect 15757 8550 15768 8676
rect 15694 8539 15768 8550
rect 1084 8370 7416 8382
rect 1084 8336 1192 8370
rect 7308 8336 7416 8370
rect 1084 8324 7416 8336
rect -27 8084 7733 8090
rect -27 8075 121 8084
rect 237 8075 7733 8084
rect -27 8041 79 8075
rect 7611 8069 7733 8075
rect 7611 8041 7649 8069
rect -27 8032 121 8041
rect 237 8032 7649 8041
rect -27 8026 7649 8032
rect -27 7979 32 8026
rect -27 79 -17 7979
rect 17 79 32 7979
rect 7643 7953 7649 8026
rect 7701 7953 7733 8069
rect 10234 8054 10292 8539
rect 15047 8452 15111 8458
rect 10953 8415 11017 8421
rect 10346 8364 10420 8375
rect 10346 8238 10357 8364
rect 10409 8238 10420 8364
rect 10953 8299 10959 8415
rect 11011 8299 11017 8415
rect 11441 8379 11505 8385
rect 10953 8293 11017 8299
rect 11254 8370 11318 8376
rect 11254 8254 11260 8370
rect 11312 8254 11318 8370
rect 11441 8263 11447 8379
rect 11499 8263 11505 8379
rect 11441 8257 11505 8263
rect 11620 8376 11684 8382
rect 11620 8260 11626 8376
rect 11678 8260 11684 8376
rect 11620 8254 11684 8260
rect 11970 8376 12034 8382
rect 11970 8260 11976 8376
rect 12028 8260 12034 8376
rect 15047 8336 15053 8452
rect 15105 8336 15111 8452
rect 15047 8330 15111 8336
rect 15305 8452 15369 8458
rect 15305 8336 15311 8452
rect 15363 8336 15369 8452
rect 15305 8330 15369 8336
rect 11970 8254 12034 8260
rect 11254 8248 11318 8254
rect 10346 8227 10420 8238
rect 10616 8192 10690 8203
rect 10616 8140 10627 8192
rect 10679 8140 10690 8192
rect 10616 8129 10690 8140
rect 10972 8192 11046 8203
rect 10972 8140 10983 8192
rect 11035 8140 11046 8192
rect 10972 8129 11046 8140
rect 11339 8202 11413 8213
rect 11339 8150 11350 8202
rect 11402 8150 11413 8202
rect 13412 8192 13540 8198
rect 11339 8139 11413 8150
rect 11747 8166 11821 8177
rect 11747 8114 11758 8166
rect 11810 8114 11821 8166
rect 13150 8140 13216 8186
rect 13412 8140 13418 8192
rect 13534 8140 13540 8192
rect 13412 8134 13540 8140
rect 13682 8191 13810 8197
rect 13682 8139 13688 8191
rect 13804 8139 13810 8191
rect 13682 8133 13810 8139
rect 14147 8187 14275 8193
rect 14147 8135 14153 8187
rect 14269 8135 14275 8187
rect 14843 8188 14971 8194
rect 14843 8186 14849 8188
rect 14522 8140 14849 8186
rect 14147 8129 14275 8135
rect 14843 8136 14849 8140
rect 14965 8136 14971 8188
rect 14843 8130 14971 8136
rect 15455 8186 15583 8192
rect 15455 8134 15461 8186
rect 15577 8134 15583 8186
rect 15455 8128 15583 8134
rect 11747 8103 11821 8114
rect 15704 8054 15762 8539
rect 10234 8042 15762 8054
rect 10234 8008 10342 8042
rect 15654 8008 15762 8042
rect 10234 7996 15762 8008
rect 7643 7947 7733 7953
rect 123 7933 251 7939
rect 123 7817 129 7933
rect 245 7817 251 7933
rect 123 7811 251 7817
rect 763 7518 879 7939
rect 1519 7518 1635 7939
rect 2275 7518 2391 7939
rect 3031 7518 3147 7939
rect 3787 7518 3903 7939
rect 4543 7518 4659 7939
rect 5299 7518 5415 7939
rect 6055 7518 6171 7939
rect 6811 7518 6927 7939
rect 7439 7933 7567 7939
rect 7439 7817 7445 7933
rect 7561 7817 7567 7933
rect 7439 7811 7567 7817
rect 7661 7911 7733 7947
rect 385 119 501 540
rect 1141 119 1257 540
rect 1897 119 2013 540
rect 2653 119 2769 540
rect 3409 119 3525 540
rect 4165 119 4281 540
rect 4921 119 5037 540
rect 5677 119 5793 540
rect 6433 119 6549 540
rect 7189 119 7305 540
rect 7661 148 7673 7911
rect 7707 148 7733 7911
rect 11908 7655 11982 7666
rect 11047 7644 11111 7650
rect 9080 7630 9144 7636
rect 9080 7578 9086 7630
rect 9138 7578 9144 7630
rect 9168 7581 10658 7627
rect 11047 7592 11053 7644
rect 11105 7592 11111 7644
rect 11047 7586 11111 7592
rect 11393 7640 11467 7651
rect 11393 7588 11404 7640
rect 11456 7588 11467 7640
rect 9080 7572 9144 7578
rect 11393 7577 11467 7588
rect 11751 7640 11825 7651
rect 11751 7588 11762 7640
rect 11814 7588 11825 7640
rect 11908 7603 11919 7655
rect 11971 7603 11982 7655
rect 11908 7592 11982 7603
rect 12533 7638 12661 7644
rect 11751 7577 11825 7588
rect 12533 7586 12539 7638
rect 12655 7586 12661 7638
rect 12533 7580 12661 7586
rect 12988 7642 13116 7648
rect 15455 7646 15583 7652
rect 12988 7590 12994 7642
rect 13110 7590 13116 7642
rect 13909 7638 14037 7644
rect 12988 7584 13116 7590
rect 13367 7581 13433 7627
rect 13909 7586 13915 7638
rect 14031 7586 14037 7638
rect 13909 7580 14037 7586
rect 14843 7636 14971 7642
rect 14843 7584 14849 7636
rect 14965 7584 14971 7636
rect 15455 7594 15461 7646
rect 15577 7594 15583 7646
rect 15455 7588 15583 7594
rect 14843 7578 14971 7584
rect 11481 7502 11545 7508
rect 10954 7494 11018 7500
rect 10954 7378 10960 7494
rect 11012 7378 11018 7494
rect 11269 7491 11333 7497
rect 11269 7467 11275 7491
rect 11182 7411 11275 7467
rect 10954 7372 11018 7378
rect 11269 7375 11275 7411
rect 11327 7375 11333 7491
rect 11481 7386 11487 7502
rect 11539 7386 11545 7502
rect 11481 7380 11545 7386
rect 11659 7502 11723 7508
rect 11659 7386 11665 7502
rect 11717 7386 11723 7502
rect 11659 7380 11723 7386
rect 12026 7502 12090 7508
rect 12026 7386 12032 7502
rect 12084 7386 12090 7502
rect 15305 7464 15369 7470
rect 12026 7380 12090 7386
rect 15043 7457 15107 7463
rect 11269 7369 11333 7375
rect 12906 7367 12980 7378
rect 9166 7335 9240 7346
rect 9166 7209 9177 7335
rect 9229 7209 9240 7335
rect 9166 7198 9240 7209
rect 9520 7335 9594 7346
rect 9520 7209 9531 7335
rect 9583 7209 9594 7335
rect 9520 7198 9594 7209
rect 9876 7335 9950 7346
rect 9876 7209 9887 7335
rect 9939 7209 9950 7335
rect 9876 7198 9950 7209
rect 10232 7335 10306 7346
rect 10232 7209 10243 7335
rect 10295 7209 10306 7335
rect 10232 7198 10306 7209
rect 10588 7335 10662 7346
rect 10588 7209 10599 7335
rect 10651 7209 10662 7335
rect 12906 7241 12917 7367
rect 12969 7241 12980 7367
rect 15043 7341 15049 7457
rect 15101 7341 15107 7457
rect 15305 7348 15311 7464
rect 15363 7348 15369 7464
rect 15305 7342 15369 7348
rect 15043 7335 15107 7341
rect 12906 7230 12980 7241
rect 10588 7198 10662 7209
rect 8984 7171 9058 7182
rect 8984 7045 8995 7171
rect 9047 7045 9058 7171
rect 8984 7034 9058 7045
rect 9342 7171 9416 7182
rect 9342 7045 9353 7171
rect 9405 7045 9416 7171
rect 9342 7034 9416 7045
rect 9698 7171 9772 7182
rect 9698 7045 9709 7171
rect 9761 7045 9772 7171
rect 9698 7034 9772 7045
rect 10054 7171 10128 7182
rect 10054 7045 10065 7171
rect 10117 7045 10128 7171
rect 10054 7034 10128 7045
rect 10410 7171 10484 7182
rect 10410 7045 10421 7171
rect 10473 7045 10484 7171
rect 10410 7034 10484 7045
rect 10766 7171 10840 7182
rect 10766 7045 10777 7171
rect 10829 7045 10840 7171
rect 10766 7034 10840 7045
rect 13812 7167 13886 7178
rect 13812 7041 13823 7167
rect 13875 7041 13886 7167
rect 13812 7030 13886 7041
rect 8852 6853 8926 6864
rect 8852 6727 8863 6853
rect 8915 6727 8926 6853
rect 8852 6716 8926 6727
rect 12146 6853 12220 6864
rect 12146 6727 12157 6853
rect 12209 6727 12220 6853
rect 12146 6716 12220 6727
rect 12314 6853 12388 6864
rect 12314 6727 12325 6853
rect 12377 6727 12388 6853
rect 12314 6716 12388 6727
rect 12447 6853 12521 6864
rect 12447 6727 12458 6853
rect 12510 6727 12521 6853
rect 12447 6716 12521 6727
rect 13363 6853 13437 6864
rect 13363 6727 13374 6853
rect 13426 6727 13437 6853
rect 13363 6716 13437 6727
rect 14279 6853 14353 6864
rect 14279 6727 14290 6853
rect 14342 6727 14353 6853
rect 14279 6716 14353 6727
rect 14413 6853 14487 6864
rect 14413 6727 14424 6853
rect 14476 6727 14487 6853
rect 14413 6716 14487 6727
rect 14654 6853 14728 6864
rect 14654 6727 14665 6853
rect 14717 6727 14728 6853
rect 14654 6716 14728 6727
rect 14788 6853 14862 6864
rect 14788 6727 14799 6853
rect 14851 6727 14862 6853
rect 14788 6716 14862 6727
rect 15562 6853 15636 6864
rect 15562 6727 15573 6853
rect 15625 6727 15636 6853
rect 15562 6716 15636 6727
rect 15696 6853 15770 6864
rect 15696 6727 15707 6853
rect 15759 6727 15770 6853
rect 15696 6716 15770 6727
rect 9080 6520 9144 6526
rect 9080 6468 9086 6520
rect 9138 6468 9144 6520
rect 10846 6522 10910 6528
rect 9168 6471 10658 6517
rect 9080 6462 9144 6468
rect 10846 6470 10852 6522
rect 10904 6470 10910 6522
rect 10846 6464 10910 6470
rect 11210 6525 11274 6531
rect 11210 6473 11216 6525
rect 11268 6473 11274 6525
rect 11210 6467 11274 6473
rect 11571 6529 11635 6535
rect 11571 6477 11577 6529
rect 11629 6477 11635 6529
rect 11571 6471 11635 6477
rect 8486 5965 15444 5977
rect 8486 5931 8594 5965
rect 15336 5931 15444 5965
rect 8486 5919 15444 5931
rect 8486 5869 8544 5919
rect 8486 5664 8498 5869
rect 8478 5653 8498 5664
rect 8532 5664 8544 5869
rect 15386 5869 15444 5919
rect 12501 5845 12629 5851
rect 8626 5787 8682 5833
rect 11932 5787 11998 5833
rect 12501 5793 12507 5845
rect 12623 5793 12629 5845
rect 12501 5787 12629 5793
rect 15248 5787 15304 5833
rect 8626 5755 8672 5787
rect 15258 5755 15304 5787
rect 15386 5664 15398 5869
rect 8532 5653 8552 5664
rect 8478 5527 8489 5653
rect 8541 5527 8552 5653
rect 8478 5516 8498 5527
rect 8486 4508 8498 5516
rect 8478 4497 8498 4508
rect 8532 5516 8552 5527
rect 8612 5653 8686 5664
rect 8612 5527 8623 5653
rect 8675 5527 8686 5653
rect 8612 5516 8686 5527
rect 10270 5653 10344 5664
rect 10270 5527 10281 5653
rect 10333 5527 10344 5653
rect 10270 5516 10344 5527
rect 13586 5653 13660 5664
rect 13586 5527 13597 5653
rect 13649 5527 13660 5653
rect 13586 5516 13660 5527
rect 15244 5653 15318 5664
rect 15244 5527 15255 5653
rect 15307 5527 15318 5653
rect 15244 5516 15318 5527
rect 15378 5653 15398 5664
rect 15432 5664 15444 5869
rect 15432 5653 15452 5664
rect 15378 5527 15389 5653
rect 15441 5527 15452 5653
rect 15378 5516 15398 5527
rect 8532 4508 8544 5516
rect 11894 5416 12042 5427
rect 11894 5364 11905 5416
rect 12031 5364 12042 5416
rect 11894 5353 11939 5364
rect 11933 5287 11939 5353
rect 11991 5353 12042 5364
rect 11991 5287 11997 5353
rect 11933 5281 11997 5287
rect 12501 4689 12629 4695
rect 8626 4631 8682 4677
rect 11932 4631 11998 4677
rect 12501 4637 12507 4689
rect 12623 4637 12629 4689
rect 12501 4631 12629 4637
rect 15248 4631 15304 4677
rect 8626 4599 8672 4631
rect 15258 4599 15304 4631
rect 15386 4508 15398 5516
rect 8532 4497 8552 4508
rect 8478 4371 8489 4497
rect 8541 4371 8552 4497
rect 8478 4360 8498 4371
rect 8486 3352 8498 4360
rect 8478 3341 8498 3352
rect 8532 4360 8552 4371
rect 8612 4497 8686 4508
rect 8612 4371 8623 4497
rect 8675 4371 8686 4497
rect 8612 4360 8686 4371
rect 10270 4497 10344 4508
rect 10270 4371 10281 4497
rect 10333 4371 10344 4497
rect 10270 4360 10344 4371
rect 13586 4497 13660 4508
rect 13586 4371 13597 4497
rect 13649 4371 13660 4497
rect 13586 4360 13660 4371
rect 15244 4497 15318 4508
rect 15244 4371 15255 4497
rect 15307 4371 15318 4497
rect 15244 4360 15318 4371
rect 15378 4497 15398 4508
rect 15432 5516 15452 5527
rect 15432 4508 15444 5516
rect 15432 4497 15452 4508
rect 15378 4371 15389 4497
rect 15441 4371 15452 4497
rect 15378 4360 15398 4371
rect 8532 3352 8544 4360
rect 11933 4247 11997 4253
rect 11933 4131 11939 4247
rect 11991 4131 11997 4247
rect 11933 4125 11997 4131
rect 12501 3533 12629 3539
rect 8626 3475 8682 3521
rect 11932 3475 11998 3521
rect 12501 3481 12507 3533
rect 12623 3481 12629 3533
rect 12501 3475 12629 3481
rect 15248 3475 15304 3521
rect 8626 3443 8672 3475
rect 11942 3443 11988 3475
rect 12542 3443 12588 3475
rect 15258 3443 15304 3475
rect 15386 3352 15398 4360
rect 8532 3341 8552 3352
rect 8478 3215 8489 3341
rect 8541 3215 8552 3341
rect 8478 3204 8498 3215
rect 8486 2196 8498 3204
rect 8478 2185 8498 2196
rect 8532 3204 8552 3215
rect 8612 3341 8686 3352
rect 8612 3215 8623 3341
rect 8675 3215 8686 3341
rect 8612 3204 8686 3215
rect 10270 3341 10344 3352
rect 10270 3215 10281 3341
rect 10333 3215 10344 3341
rect 10270 3204 10344 3215
rect 13586 3341 13660 3352
rect 13586 3215 13597 3341
rect 13649 3215 13660 3341
rect 13586 3204 13660 3215
rect 15244 3341 15318 3352
rect 15244 3215 15255 3341
rect 15307 3215 15318 3341
rect 15244 3204 15318 3215
rect 15378 3341 15398 3352
rect 15432 4360 15452 4371
rect 15432 3352 15444 4360
rect 15432 3341 15452 3352
rect 15378 3215 15389 3341
rect 15441 3215 15452 3341
rect 15378 3204 15398 3215
rect 8532 2196 8544 3204
rect 11674 2998 11738 3004
rect 11674 2882 11680 2998
rect 11732 2968 11738 2998
rect 11732 2914 11954 2968
rect 11732 2882 11738 2914
rect 11674 2876 11738 2882
rect 12501 2377 12629 2383
rect 8626 2319 8682 2365
rect 11932 2319 11998 2365
rect 12501 2325 12507 2377
rect 12623 2325 12629 2377
rect 12501 2319 12629 2325
rect 15248 2319 15304 2365
rect 8626 2287 8672 2319
rect 15258 2287 15304 2319
rect 15386 2196 15398 3204
rect 8532 2185 8552 2196
rect 8478 2059 8489 2185
rect 8541 2059 8552 2185
rect 8478 2048 8498 2059
rect 8486 1040 8498 2048
rect 8478 1029 8498 1040
rect 8532 2048 8552 2059
rect 8612 2185 8686 2196
rect 8612 2059 8623 2185
rect 8675 2059 8686 2185
rect 8612 2048 8686 2059
rect 10270 2185 10344 2196
rect 10270 2059 10281 2185
rect 10333 2059 10344 2185
rect 10270 2048 10344 2059
rect 13586 2185 13660 2196
rect 13586 2059 13597 2185
rect 13649 2059 13660 2185
rect 13586 2048 13660 2059
rect 15244 2185 15318 2196
rect 15244 2059 15255 2185
rect 15307 2059 15318 2185
rect 15244 2048 15318 2059
rect 15378 2185 15398 2196
rect 15432 3204 15452 3215
rect 15432 2196 15444 3204
rect 15432 2185 15452 2196
rect 15378 2059 15389 2185
rect 15441 2059 15452 2185
rect 15378 2048 15398 2059
rect 8532 1040 8544 2048
rect 11933 1935 11997 1941
rect 11933 1819 11939 1935
rect 11991 1819 11997 1935
rect 11933 1813 11997 1819
rect 12501 1221 12629 1227
rect 8626 1163 8682 1209
rect 11932 1163 11998 1209
rect 12501 1169 12507 1221
rect 12623 1169 12629 1221
rect 12501 1163 12629 1169
rect 15248 1163 15304 1209
rect 8626 1131 8672 1163
rect 15258 1131 15304 1163
rect 15386 1040 15398 2048
rect 8532 1029 8552 1040
rect 8478 903 8489 1029
rect 8541 903 8552 1029
rect 8478 892 8498 903
rect 7661 138 7733 148
rect 7660 111 7733 138
rect -27 33 32 79
rect 7643 105 7733 111
rect 7643 33 7649 105
rect -27 17 7649 33
rect -27 -17 79 17
rect 7611 -11 7649 17
rect 7701 -11 7733 105
rect 7611 -17 7733 -11
rect -27 -27 7733 -17
rect 8486 79 8498 892
rect 8532 892 8552 903
rect 8612 1029 8686 1040
rect 8612 903 8623 1029
rect 8675 903 8686 1029
rect 8612 892 8686 903
rect 10270 1029 10344 1040
rect 10270 903 10281 1029
rect 10333 903 10344 1029
rect 10270 892 10344 903
rect 13586 1029 13660 1040
rect 13586 903 13597 1029
rect 13649 903 13660 1029
rect 13586 892 13660 903
rect 15244 1029 15318 1040
rect 15244 903 15255 1029
rect 15307 903 15318 1029
rect 15244 892 15318 903
rect 15378 1029 15398 1040
rect 15432 2048 15452 2059
rect 15432 1040 15444 2048
rect 15432 1029 15452 1040
rect 15378 903 15389 1029
rect 15441 903 15452 1029
rect 15378 892 15398 903
rect 8532 79 8544 892
rect 11933 779 11997 785
rect 11933 663 11939 779
rect 11991 663 11997 779
rect 11933 657 11997 663
rect 8486 29 8544 79
rect 15386 79 15398 892
rect 15432 892 15452 903
rect 15432 79 15444 892
rect 15386 29 15444 79
rect 8486 17 15444 29
rect 8486 -17 8594 17
rect 15336 -17 15444 17
rect -27 -63 32 -27
rect 8486 -29 15444 -17
rect -138 -69 8047 -63
rect -138 -346 7751 -69
rect 8041 -346 8047 -69
rect -138 -352 8047 -346
rect -138 -408 8402 -402
rect -138 -646 8106 -408
rect 8396 -646 8402 -408
rect -138 -652 8402 -646
<< via1 >>
rect 3651 11255 3777 11307
rect 4723 11255 4849 11307
rect 8085 11066 8137 11192
rect 9801 11066 9853 11192
rect 1084 10697 1136 10711
rect 1084 10599 1093 10697
rect 1093 10599 1127 10697
rect 1127 10599 1136 10697
rect 1084 10585 1136 10599
rect 1220 10585 1272 10711
rect 2078 10585 2130 10711
rect 3794 10585 3846 10711
rect 4652 10585 4704 10711
rect 6368 10585 6420 10711
rect 7227 10585 7279 10711
rect 8943 10585 8995 10711
rect 10659 10585 10711 10711
rect 12375 10585 12427 10711
rect 13233 10585 13285 10711
rect 13366 10697 13418 10711
rect 13366 10599 13375 10697
rect 13375 10599 13409 10697
rect 13409 10599 13418 10697
rect 13366 10585 13418 10599
rect 2937 10209 2989 10325
rect 5511 10209 5563 10325
rect 3651 10099 3777 10151
rect 4723 10099 4849 10151
rect 10261 10120 10377 10172
rect 11433 10131 11549 10183
rect 3651 9595 3777 9647
rect 4723 9595 4849 9647
rect 2937 9430 2989 9546
rect 5511 9430 5563 9546
rect 1084 9197 1136 9211
rect 1084 9099 1093 9197
rect 1093 9099 1127 9197
rect 1127 9099 1136 9197
rect 1084 9085 1136 9099
rect 1220 9085 1272 9211
rect 4227 9085 4279 9137
rect 2079 8634 2131 8760
rect 3795 8634 3847 8760
rect 7227 9085 7279 9211
rect 7361 9197 7413 9211
rect 7361 9099 7370 9197
rect 7370 9099 7404 9197
rect 7404 9099 7413 9197
rect 7361 9085 7413 9099
rect 4653 8634 4705 8760
rect 6369 8634 6421 8760
rect 3651 8445 3777 8497
rect 4723 8445 4849 8497
rect 10464 9275 10516 9327
rect 10618 9270 10670 9322
rect 10825 9257 10877 9309
rect 11172 9265 11224 9317
rect 11528 9265 11580 9317
rect 11882 9266 11934 9318
rect 12326 9270 12442 9322
rect 10943 9014 10995 9140
rect 13616 9053 13668 9179
rect 11048 8792 11100 8918
rect 12695 8884 12747 9010
rect 14534 8768 14586 8894
rect 10237 8662 10289 8676
rect 10237 8564 10246 8662
rect 10246 8564 10280 8662
rect 10280 8564 10289 8662
rect 10237 8550 10289 8564
rect 10727 8655 10779 8707
rect 12105 8662 12157 8676
rect 12105 8564 12114 8662
rect 12114 8564 12148 8662
rect 12148 8564 12157 8662
rect 12105 8550 12157 8564
rect 12241 8550 12293 8676
rect 13157 8550 13209 8676
rect 14073 8550 14125 8676
rect 14665 8662 14717 8676
rect 14665 8564 14674 8662
rect 14674 8564 14708 8662
rect 14708 8564 14717 8662
rect 14665 8550 14717 8564
rect 14799 8550 14851 8676
rect 15573 8550 15625 8676
rect 15705 8550 15757 8676
rect 121 8075 237 8084
rect 121 8041 237 8075
rect 7649 8060 7701 8069
rect 121 8032 237 8041
rect 7649 7962 7658 8060
rect 7658 7962 7692 8060
rect 7692 7962 7701 8060
rect 7649 7953 7701 7962
rect 10357 8238 10409 8364
rect 10959 8299 11011 8415
rect 11260 8254 11312 8370
rect 11447 8263 11499 8379
rect 11626 8260 11678 8376
rect 11976 8260 12028 8376
rect 15053 8336 15105 8452
rect 15311 8336 15363 8452
rect 10627 8140 10679 8192
rect 10983 8140 11035 8192
rect 11350 8150 11402 8202
rect 11758 8114 11810 8166
rect 13418 8140 13534 8192
rect 13688 8139 13804 8191
rect 14153 8135 14269 8187
rect 14849 8136 14965 8188
rect 15461 8134 15577 8186
rect 129 7817 245 7933
rect 7445 7817 7561 7933
rect 9086 7578 9138 7630
rect 11053 7592 11105 7644
rect 11404 7588 11456 7640
rect 11762 7588 11814 7640
rect 11919 7603 11971 7655
rect 12539 7586 12655 7638
rect 12994 7590 13110 7642
rect 13915 7586 14031 7638
rect 14849 7584 14965 7636
rect 15461 7594 15577 7646
rect 10960 7378 11012 7494
rect 11275 7375 11327 7491
rect 11487 7386 11539 7502
rect 11665 7386 11717 7502
rect 12032 7386 12084 7502
rect 9177 7209 9229 7335
rect 9531 7209 9583 7335
rect 9887 7209 9939 7335
rect 10243 7209 10295 7335
rect 10599 7209 10651 7335
rect 12917 7241 12969 7367
rect 15049 7341 15101 7457
rect 15311 7348 15363 7464
rect 8995 7045 9047 7171
rect 9353 7045 9405 7171
rect 9709 7045 9761 7171
rect 10065 7045 10117 7171
rect 10421 7045 10473 7171
rect 10777 7045 10829 7171
rect 13823 7041 13875 7167
rect 8863 6839 8915 6853
rect 8863 6741 8872 6839
rect 8872 6741 8906 6839
rect 8906 6741 8915 6839
rect 8863 6727 8915 6741
rect 12157 6839 12209 6853
rect 12157 6741 12166 6839
rect 12166 6741 12200 6839
rect 12200 6741 12209 6839
rect 12157 6727 12209 6741
rect 12325 6839 12377 6853
rect 12325 6741 12334 6839
rect 12334 6741 12368 6839
rect 12368 6741 12377 6839
rect 12325 6727 12377 6741
rect 12458 6727 12510 6853
rect 13374 6727 13426 6853
rect 14290 6727 14342 6853
rect 14424 6839 14476 6853
rect 14424 6741 14433 6839
rect 14433 6741 14467 6839
rect 14467 6741 14476 6839
rect 14424 6727 14476 6741
rect 14665 6727 14717 6853
rect 14799 6727 14851 6853
rect 15573 6727 15625 6853
rect 15707 6727 15759 6853
rect 9086 6468 9138 6520
rect 10852 6470 10904 6522
rect 11216 6473 11268 6525
rect 11577 6477 11629 6529
rect 12507 5793 12623 5845
rect 8489 5527 8498 5653
rect 8498 5527 8532 5653
rect 8532 5527 8541 5653
rect 8623 5527 8675 5653
rect 10281 5527 10333 5653
rect 13597 5527 13649 5653
rect 15255 5527 15307 5653
rect 15389 5527 15398 5653
rect 15398 5527 15432 5653
rect 15432 5527 15441 5653
rect 11905 5364 12031 5416
rect 11939 5287 11991 5364
rect 12507 4637 12623 4689
rect 8489 4371 8498 4497
rect 8498 4371 8532 4497
rect 8532 4371 8541 4497
rect 8623 4371 8675 4497
rect 10281 4371 10333 4497
rect 13597 4371 13649 4497
rect 15255 4371 15307 4497
rect 15389 4371 15398 4497
rect 15398 4371 15432 4497
rect 15432 4371 15441 4497
rect 11939 4131 11991 4247
rect 12507 3481 12623 3533
rect 8489 3215 8498 3341
rect 8498 3215 8532 3341
rect 8532 3215 8541 3341
rect 8623 3215 8675 3341
rect 10281 3215 10333 3341
rect 13597 3215 13649 3341
rect 15255 3215 15307 3341
rect 15389 3215 15398 3341
rect 15398 3215 15432 3341
rect 15432 3215 15441 3341
rect 11680 2882 11732 2998
rect 12507 2325 12623 2377
rect 8489 2059 8498 2185
rect 8498 2059 8532 2185
rect 8532 2059 8541 2185
rect 8623 2059 8675 2185
rect 10281 2059 10333 2185
rect 13597 2059 13649 2185
rect 15255 2059 15307 2185
rect 15389 2059 15398 2185
rect 15398 2059 15432 2185
rect 15432 2059 15441 2185
rect 11939 1819 11991 1935
rect 12507 1169 12623 1221
rect 8489 903 8498 1029
rect 8498 903 8532 1029
rect 8532 903 8541 1029
rect 7649 96 7701 105
rect 7649 -2 7658 96
rect 7658 -2 7692 96
rect 7692 -2 7701 96
rect 7649 -11 7701 -2
rect 8623 903 8675 1029
rect 10281 903 10333 1029
rect 13597 903 13649 1029
rect 15255 903 15307 1029
rect 15389 903 15398 1029
rect 15398 903 15432 1029
rect 15432 903 15441 1029
rect 11939 663 11991 779
rect 7751 -346 8041 -69
rect 8106 -646 8396 -408
<< metal2 >>
rect 3640 11309 3788 11318
rect 3640 11253 3649 11309
rect 3779 11253 3788 11309
rect 3640 11244 3788 11253
rect 4712 11309 4860 11318
rect 4712 11253 4721 11309
rect 4851 11253 4860 11309
rect 4712 11244 4860 11253
rect 8074 11194 8148 11203
rect 8074 11064 8083 11194
rect 8139 11064 8148 11194
rect 8074 11055 8148 11064
rect 9790 11194 9864 11203
rect 9790 11064 9799 11194
rect 9855 11064 9864 11194
rect 9790 11055 9864 11064
rect 1073 10713 1147 10722
rect 1073 10583 1082 10713
rect 1138 10583 1147 10713
rect 1073 10574 1147 10583
rect 1209 10713 1283 10722
rect 1209 10583 1218 10713
rect 1274 10583 1283 10713
rect 1209 10574 1283 10583
rect 2067 10713 2141 10722
rect 2067 10583 2076 10713
rect 2132 10583 2141 10713
rect 2067 10574 2141 10583
rect 3783 10713 3857 10722
rect 3783 10583 3792 10713
rect 3848 10583 3857 10713
rect 3783 10574 3857 10583
rect 4641 10713 4715 10722
rect 4641 10583 4650 10713
rect 4706 10583 4715 10713
rect 4641 10574 4715 10583
rect 6357 10713 6431 10722
rect 6357 10583 6366 10713
rect 6422 10583 6431 10713
rect 6357 10574 6431 10583
rect 7216 10713 7290 10722
rect 7216 10583 7225 10713
rect 7281 10583 7290 10713
rect 7216 10574 7290 10583
rect 8100 10709 8402 10721
rect 8100 10589 8113 10709
rect 8382 10589 8402 10709
rect 2931 10325 2995 10331
rect 2931 10209 2937 10325
rect 2989 10209 2995 10325
rect 2931 9546 2995 10209
rect 5505 10325 5569 10331
rect 5505 10209 5511 10325
rect 5563 10209 5569 10325
rect 3640 10153 3788 10162
rect 3640 10097 3649 10153
rect 3779 10097 3788 10153
rect 3640 10088 3788 10097
rect 4712 10153 4860 10162
rect 4712 10097 4721 10153
rect 4851 10097 4860 10153
rect 4712 10088 4860 10097
rect 3640 9649 3788 9658
rect 3640 9593 3649 9649
rect 3779 9593 3788 9649
rect 3640 9584 3788 9593
rect 4712 9649 4860 9658
rect 4712 9593 4721 9649
rect 4851 9593 4860 9649
rect 4712 9584 4860 9593
rect 2931 9430 2937 9546
rect 2989 9430 2995 9546
rect 2931 9424 2995 9430
rect 5505 9546 5569 10209
rect 5505 9430 5511 9546
rect 5563 9430 5569 9546
rect 5505 9428 5569 9430
rect 5504 9424 5569 9428
rect 141 9213 215 9222
rect 141 9083 150 9213
rect 206 9083 215 9213
rect 141 9074 215 9083
rect 1073 9213 1147 9222
rect 1073 9083 1082 9213
rect 1138 9083 1147 9213
rect 1073 9074 1147 9083
rect 1209 9213 1283 9222
rect 1209 9083 1218 9213
rect 1274 9083 1283 9213
rect 1209 9074 1283 9083
rect 4216 9139 4290 9148
rect 4216 9083 4225 9139
rect 4281 9083 4290 9139
rect 4216 9074 4290 9083
rect 147 8090 211 9074
rect 2068 8762 2142 8771
rect 2068 8632 2077 8762
rect 2133 8632 2142 8762
rect 2068 8623 2142 8632
rect 3784 8762 3858 8771
rect 3784 8632 3793 8762
rect 3849 8632 3858 8762
rect 3784 8623 3858 8632
rect 4642 8762 4716 8771
rect 4642 8632 4651 8762
rect 4707 8632 4716 8762
rect 4642 8623 4716 8632
rect 3640 8499 3788 8508
rect 3640 8443 3649 8499
rect 3779 8443 3788 8499
rect 3640 8434 3788 8443
rect 4712 8499 4860 8508
rect 4712 8443 4721 8499
rect 4851 8443 4860 8499
rect 4712 8434 4860 8443
rect 115 8084 243 8090
rect 115 8032 121 8084
rect 237 8032 243 8084
rect 5504 8065 5566 9424
rect 7216 9213 7290 9222
rect 7216 9083 7225 9213
rect 7281 9083 7290 9213
rect 7216 9074 7290 9083
rect 7350 9213 7424 9222
rect 7350 9083 7359 9213
rect 7415 9083 7424 9213
rect 7350 9074 7424 9083
rect 7745 9213 8047 9790
rect 7745 9083 7754 9213
rect 7810 9083 8047 9213
rect 6358 8762 6432 8771
rect 6358 8632 6367 8762
rect 6423 8632 6432 8762
rect 6358 8623 6432 8632
rect 7430 8739 7504 8748
rect 7430 8609 7439 8739
rect 7495 8609 7504 8739
rect 7430 8600 7504 8609
rect 6934 8521 7008 8530
rect 6934 8391 6943 8521
rect 6999 8391 7008 8521
rect 6934 8382 7008 8391
rect 115 8026 243 8032
rect 5498 8056 5572 8065
rect 147 7939 211 8026
rect 123 7933 251 7939
rect 123 7817 129 7933
rect 245 7817 251 7933
rect 5498 7926 5507 8056
rect 5563 7926 5572 8056
rect 5498 7917 5572 7926
rect 123 7811 251 7817
rect 6946 7157 7008 8382
rect 7444 7939 7500 8600
rect 7745 8075 8047 9083
rect 7643 8069 8047 8075
rect 7643 7953 7649 8069
rect 7701 7953 8047 8069
rect 7643 7947 8047 7953
rect 7439 7933 7567 7939
rect 7439 7817 7445 7933
rect 7561 7817 7567 7933
rect 7439 7811 7567 7817
rect 6942 7148 7016 7157
rect 6942 7018 6951 7148
rect 7007 7018 7016 7148
rect 6942 7009 7016 7018
rect 7745 6855 8047 7947
rect 7745 6725 7982 6855
rect 8038 6725 8047 6855
rect 7745 5655 8047 6725
rect 7745 5525 7982 5655
rect 8038 5525 8047 5655
rect 7745 4499 8047 5525
rect 7745 4369 7982 4499
rect 8038 4369 8047 4499
rect 7745 3343 8047 4369
rect 7745 3213 7982 3343
rect 8038 3213 8047 3343
rect 7745 2187 8047 3213
rect 7745 2057 7982 2187
rect 8038 2057 8047 2187
rect 7745 1031 8047 2057
rect 7745 901 7982 1031
rect 8038 901 8047 1031
rect 7745 111 8047 901
rect 7643 105 8047 111
rect 7643 -11 7649 105
rect 7701 -11 8047 105
rect 7643 -17 8047 -11
rect 7745 -69 8047 -17
rect 7745 -346 7751 -69
rect 8041 -346 8047 -69
rect 7745 -352 8047 -346
rect 8100 8678 8402 10589
rect 8932 10713 9006 10722
rect 8932 10583 8941 10713
rect 8997 10583 9006 10713
rect 8932 10574 9006 10583
rect 10648 10713 10722 10722
rect 10648 10583 10657 10713
rect 10713 10583 10722 10713
rect 10648 10574 10722 10583
rect 12364 10713 12438 10722
rect 12364 10583 12373 10713
rect 12429 10583 12438 10713
rect 12364 10574 12438 10583
rect 13222 10713 13296 10722
rect 13222 10583 13231 10713
rect 13287 10583 13296 10713
rect 13222 10574 13296 10583
rect 13355 10713 13429 10722
rect 13355 10583 13364 10713
rect 13420 10583 13429 10713
rect 13355 10574 13429 10583
rect 11427 10183 11555 10189
rect 10255 10172 10383 10178
rect 10255 10120 10261 10172
rect 10377 10120 10383 10172
rect 11427 10131 11433 10183
rect 11549 10131 11555 10183
rect 11427 10125 11555 10131
rect 10255 10114 10383 10120
rect 10288 9007 10356 10114
rect 10601 9547 10749 9556
rect 10601 9491 10610 9547
rect 10740 9491 10749 9547
rect 10601 9482 10749 9491
rect 10453 9329 10527 9338
rect 10453 9273 10462 9329
rect 10518 9273 10527 9329
rect 10453 9264 10527 9273
rect 10609 9322 10678 9482
rect 10609 9270 10618 9322
rect 10670 9270 10678 9322
rect 11166 9317 11230 9323
rect 10276 8998 10356 9007
rect 10276 8868 10285 8998
rect 10341 8868 10356 8998
rect 10276 8860 10356 8868
rect 10276 8859 10350 8860
rect 8100 8548 8337 8678
rect 8393 8548 8402 8678
rect 8100 -408 8402 8548
rect 10226 8678 10300 8687
rect 10226 8548 10235 8678
rect 10291 8548 10300 8678
rect 10226 8539 10300 8548
rect 10346 8366 10420 8375
rect 10346 8236 10355 8366
rect 10411 8236 10420 8366
rect 10346 8227 10420 8236
rect 9080 7630 9144 7636
rect 9080 7578 9086 7630
rect 9138 7578 9144 7630
rect 9080 7572 9144 7578
rect 8984 7173 9058 7182
rect 8984 7043 8993 7173
rect 9049 7043 9058 7173
rect 8984 7034 9058 7043
rect 8852 6855 8926 6864
rect 8852 6725 8861 6855
rect 8917 6725 8926 6855
rect 8852 6716 8926 6725
rect 9086 6526 9138 7572
rect 10346 7529 10400 8227
rect 10609 8203 10678 9270
rect 10819 9309 10883 9315
rect 10819 9257 10825 9309
rect 10877 9257 10883 9309
rect 10716 8709 10790 8718
rect 10716 8653 10725 8709
rect 10781 8653 10790 8709
rect 10716 8644 10790 8653
rect 10819 8614 10883 9257
rect 11166 9265 11172 9317
rect 11224 9265 11230 9317
rect 10932 9142 11006 9151
rect 10932 9012 10941 9142
rect 10997 9012 11006 9142
rect 10932 9003 11006 9012
rect 11037 8920 11111 8929
rect 11037 8790 11046 8920
rect 11102 8790 11111 8920
rect 11037 8781 11111 8790
rect 11166 8614 11230 9265
rect 11435 9029 11491 10125
rect 12295 9543 12443 9552
rect 12295 9487 12304 9543
rect 12434 9487 12443 9543
rect 12295 9478 12443 9487
rect 13893 9545 14041 9554
rect 13893 9489 13902 9545
rect 14032 9489 14041 9545
rect 13893 9480 14041 9489
rect 15402 9545 15550 9554
rect 15402 9489 15411 9545
rect 15541 9489 15550 9545
rect 15402 9480 15550 9489
rect 11417 9020 11491 9029
rect 11417 8890 11426 9020
rect 11482 8890 11491 9020
rect 11417 8881 11491 8890
rect 11435 8642 11491 8881
rect 11522 9317 11586 9323
rect 11522 9265 11528 9317
rect 11580 9265 11586 9317
rect 10805 8606 10883 8614
rect 10805 8605 10879 8606
rect 10805 8549 10814 8605
rect 10870 8549 10879 8605
rect 10805 8540 10879 8549
rect 11161 8605 11235 8614
rect 11161 8549 11170 8605
rect 11226 8549 11235 8605
rect 11161 8540 11235 8549
rect 11435 8512 11489 8642
rect 11522 8614 11586 9265
rect 11871 9320 11945 9329
rect 12345 9328 12409 9478
rect 11871 9264 11880 9320
rect 11936 9264 11945 9320
rect 12320 9322 12448 9328
rect 12320 9270 12326 9322
rect 12442 9270 12448 9322
rect 12320 9264 12448 9270
rect 11871 9255 11945 9264
rect 11517 8605 11591 8614
rect 11517 8549 11526 8605
rect 11582 8549 11591 8605
rect 11517 8540 11591 8549
rect 10953 8415 11017 8421
rect 10953 8355 10959 8415
rect 10875 8299 10959 8355
rect 11011 8299 11017 8415
rect 11435 8385 11491 8512
rect 11435 8379 11505 8385
rect 11254 8370 11318 8376
rect 11254 8328 11260 8370
rect 10875 8293 11017 8299
rect 10609 8202 10690 8203
rect 10616 8194 10690 8202
rect 10616 8138 10625 8194
rect 10681 8138 10690 8194
rect 10616 8129 10690 8138
rect 10875 8037 10931 8293
rect 11242 8254 11260 8328
rect 11312 8254 11318 8370
rect 11435 8349 11447 8379
rect 11441 8263 11447 8349
rect 11499 8306 11505 8379
rect 11620 8376 11684 8382
rect 11499 8263 11552 8306
rect 11441 8257 11552 8263
rect 11242 8248 11318 8254
rect 10972 8194 11046 8203
rect 10972 8138 10981 8194
rect 11037 8176 11046 8194
rect 11037 8138 11088 8176
rect 10972 8129 11088 8138
rect 11029 8053 11088 8129
rect 11029 8044 11104 8053
rect 10875 8001 10977 8037
rect 10875 7961 10896 8001
rect 10887 7945 10896 7961
rect 10952 7945 10977 8001
rect 11029 7988 11039 8044
rect 11095 7988 11104 8044
rect 11029 7979 11104 7988
rect 10887 7936 10977 7945
rect 10337 7520 10411 7529
rect 10337 7390 10346 7520
rect 10402 7390 10411 7520
rect 10919 7500 10977 7936
rect 11039 7902 11113 7911
rect 11039 7846 11048 7902
rect 11104 7846 11113 7902
rect 11039 7837 11113 7846
rect 11048 7650 11105 7837
rect 11047 7644 11111 7650
rect 11047 7592 11053 7644
rect 11105 7592 11111 7644
rect 11047 7586 11111 7592
rect 10919 7494 11018 7500
rect 10919 7450 10960 7494
rect 10337 7381 10411 7390
rect 10954 7378 10960 7450
rect 11012 7378 11018 7494
rect 11242 7497 11294 8248
rect 11339 8204 11413 8213
rect 11339 8148 11348 8204
rect 11404 8148 11413 8204
rect 11339 8139 11413 8148
rect 11496 8183 11552 8257
rect 11620 8260 11626 8376
rect 11678 8317 11684 8376
rect 11678 8260 11691 8317
rect 11620 8254 11691 8260
rect 11496 8146 11578 8183
rect 11343 7913 11403 8139
rect 11336 7904 11410 7913
rect 11336 7848 11345 7904
rect 11401 7848 11410 7904
rect 11336 7839 11410 7848
rect 11393 7642 11467 7651
rect 11393 7586 11402 7642
rect 11458 7586 11467 7642
rect 11393 7577 11467 7586
rect 11517 7508 11578 8146
rect 11635 8028 11691 8254
rect 11874 8212 11930 9255
rect 13605 9181 13679 9190
rect 13605 9051 13614 9181
rect 13670 9051 13679 9181
rect 13605 9042 13679 9051
rect 12684 9012 12758 9021
rect 12684 8882 12693 9012
rect 12749 8882 12758 9012
rect 12684 8873 12758 8882
rect 12094 8678 12168 8687
rect 12094 8548 12103 8678
rect 12159 8548 12168 8678
rect 12094 8539 12168 8548
rect 12230 8678 12304 8687
rect 12230 8548 12239 8678
rect 12295 8548 12304 8678
rect 12230 8539 12304 8548
rect 13146 8678 13220 8687
rect 13146 8548 13155 8678
rect 13211 8548 13220 8678
rect 13146 8539 13220 8548
rect 11970 8376 12034 8382
rect 11970 8260 11976 8376
rect 12028 8311 12034 8376
rect 12028 8260 12090 8311
rect 11970 8254 12090 8260
rect 11747 8168 11821 8177
rect 11747 8112 11756 8168
rect 11812 8112 11821 8168
rect 11874 8164 11964 8212
rect 11747 8103 11821 8112
rect 11908 8042 11964 8164
rect 11779 8032 11853 8041
rect 11635 7981 11723 8028
rect 11779 7984 11788 8032
rect 11481 7502 11578 7508
rect 11242 7491 11333 7497
rect 11242 7435 11275 7491
rect 10954 7372 11018 7378
rect 11269 7375 11275 7435
rect 11327 7375 11333 7491
rect 11481 7400 11487 7502
rect 11269 7369 11333 7375
rect 11468 7386 11487 7400
rect 11539 7475 11578 7502
rect 11659 7502 11723 7981
rect 11772 7976 11788 7984
rect 11844 7976 11853 8032
rect 11772 7967 11853 7976
rect 11908 8033 11998 8042
rect 11908 7977 11933 8033
rect 11989 7977 11998 8033
rect 11908 7968 11998 7977
rect 11772 7651 11830 7967
rect 11751 7642 11830 7651
rect 11751 7586 11760 7642
rect 11816 7636 11830 7642
rect 11908 7657 11982 7666
rect 11816 7586 11825 7636
rect 11908 7601 11917 7657
rect 11973 7601 11982 7657
rect 11908 7592 11982 7601
rect 11751 7577 11825 7586
rect 11539 7386 11545 7475
rect 11468 7380 11545 7386
rect 11659 7386 11665 7502
rect 11717 7401 11723 7502
rect 12026 7502 12090 8254
rect 13412 8192 13540 8198
rect 13412 8140 13418 8192
rect 13534 8140 13540 8192
rect 13412 8134 13540 8140
rect 13682 8191 13810 8197
rect 13682 8139 13688 8191
rect 13804 8139 13810 8191
rect 12973 8036 13121 8045
rect 12973 7980 12982 8036
rect 13112 7980 13121 8036
rect 12973 7971 13121 7980
rect 12552 7902 12626 7911
rect 12552 7846 12561 7902
rect 12617 7846 12626 7902
rect 12552 7837 12626 7846
rect 12560 7644 12617 7837
rect 13032 7648 13088 7971
rect 13460 7736 13518 8134
rect 13682 8133 13810 8139
rect 13705 7915 13766 8133
rect 13698 7906 13772 7915
rect 13698 7850 13707 7906
rect 13763 7850 13772 7906
rect 13698 7841 13772 7850
rect 13452 7727 13526 7736
rect 13452 7671 13461 7727
rect 13517 7671 13526 7727
rect 13452 7662 13526 7671
rect 12533 7638 12661 7644
rect 12533 7586 12539 7638
rect 12655 7586 12661 7638
rect 12533 7580 12661 7586
rect 12988 7642 13116 7648
rect 13936 7644 13993 9480
rect 14523 8896 14597 8905
rect 14523 8766 14532 8896
rect 14588 8766 14597 8896
rect 14523 8757 14597 8766
rect 14062 8678 14136 8687
rect 14062 8548 14071 8678
rect 14127 8548 14136 8678
rect 14062 8539 14136 8548
rect 14654 8678 14728 8687
rect 14654 8548 14663 8678
rect 14719 8548 14728 8678
rect 14654 8539 14728 8548
rect 14788 8678 14862 8687
rect 14788 8548 14797 8678
rect 14853 8548 14862 8678
rect 14788 8539 14862 8548
rect 15047 8452 15111 8458
rect 15047 8336 15053 8452
rect 15105 8389 15111 8452
rect 15305 8452 15369 8458
rect 15305 8393 15311 8452
rect 15105 8336 15139 8389
rect 15047 8330 15139 8336
rect 14147 8187 14275 8193
rect 14147 8135 14153 8187
rect 14269 8135 14275 8187
rect 14147 8129 14275 8135
rect 14843 8188 14971 8194
rect 14843 8136 14849 8188
rect 14965 8136 14971 8188
rect 14843 8130 14971 8136
rect 14165 7741 14237 8129
rect 14165 7732 14241 7741
rect 14165 7722 14176 7732
rect 14167 7676 14176 7722
rect 14232 7676 14241 7732
rect 14167 7667 14241 7676
rect 12988 7590 12994 7642
rect 13110 7590 13116 7642
rect 12988 7584 13116 7590
rect 13909 7638 14037 7644
rect 14879 7642 14933 8130
rect 15083 8038 15139 8330
rect 15267 8336 15311 8393
rect 15363 8336 15369 8452
rect 15267 8330 15369 8336
rect 15072 8029 15146 8038
rect 15072 7973 15081 8029
rect 15137 7973 15146 8029
rect 15072 7964 15146 7973
rect 13909 7586 13915 7638
rect 14031 7586 14037 7638
rect 13909 7580 14037 7586
rect 14843 7636 14971 7642
rect 14843 7584 14849 7636
rect 14965 7584 14971 7636
rect 14843 7578 14971 7584
rect 11717 7386 11732 7401
rect 11659 7380 11732 7386
rect 12026 7386 12032 7502
rect 12084 7386 12090 7502
rect 15083 7463 15139 7964
rect 15267 7908 15323 8330
rect 15470 8192 15526 9480
rect 15562 8678 15636 8687
rect 15562 8548 15571 8678
rect 15627 8548 15636 8678
rect 15562 8539 15636 8548
rect 15694 8678 15768 8687
rect 15694 8548 15703 8678
rect 15759 8548 15768 8678
rect 15694 8539 15768 8548
rect 15455 8186 15583 8192
rect 15455 8134 15461 8186
rect 15577 8134 15583 8186
rect 15455 8128 15583 8134
rect 15257 7899 15331 7908
rect 15257 7843 15266 7899
rect 15322 7843 15331 7899
rect 15257 7834 15331 7843
rect 12026 7380 12090 7386
rect 15043 7457 15139 7463
rect 9166 7337 9240 7346
rect 9166 7207 9175 7337
rect 9231 7207 9240 7337
rect 9166 7198 9240 7207
rect 9520 7337 9594 7346
rect 9520 7207 9529 7337
rect 9585 7207 9594 7337
rect 9520 7198 9594 7207
rect 9876 7337 9950 7346
rect 9876 7207 9885 7337
rect 9941 7207 9950 7337
rect 9876 7198 9950 7207
rect 10232 7337 10306 7346
rect 10232 7207 10241 7337
rect 10297 7207 10306 7337
rect 10232 7198 10306 7207
rect 10588 7337 10662 7346
rect 10588 7207 10597 7337
rect 10653 7207 10662 7337
rect 10588 7198 10662 7207
rect 9342 7173 9416 7182
rect 9342 7043 9351 7173
rect 9407 7043 9416 7173
rect 9342 7034 9416 7043
rect 9698 7173 9772 7182
rect 9698 7043 9707 7173
rect 9763 7043 9772 7173
rect 9698 7034 9772 7043
rect 10054 7173 10128 7182
rect 10054 7043 10063 7173
rect 10119 7043 10128 7173
rect 10054 7034 10128 7043
rect 10410 7173 10484 7182
rect 10410 7043 10419 7173
rect 10475 7043 10484 7173
rect 10410 7034 10484 7043
rect 10766 7173 10840 7182
rect 10766 7043 10775 7173
rect 10831 7043 10840 7173
rect 10766 7034 10840 7043
rect 10851 6793 10925 6802
rect 10851 6737 10860 6793
rect 10916 6737 10925 6793
rect 10851 6728 10925 6737
rect 11207 6794 11281 6803
rect 11207 6738 11216 6794
rect 11272 6738 11281 6794
rect 11207 6729 11281 6738
rect 10857 6528 10909 6728
rect 11213 6531 11272 6729
rect 9080 6520 9144 6526
rect 9080 6468 9086 6520
rect 9138 6468 9144 6520
rect 9080 6462 9144 6468
rect 10846 6522 10910 6528
rect 10846 6470 10852 6522
rect 10904 6470 10910 6522
rect 10846 6464 10910 6470
rect 11210 6525 11274 6531
rect 11210 6473 11216 6525
rect 11268 6473 11274 6525
rect 11210 6467 11274 6473
rect 8478 5655 8552 5664
rect 8478 5525 8487 5655
rect 8543 5525 8552 5655
rect 8478 5516 8552 5525
rect 8612 5655 8686 5664
rect 8612 5525 8621 5655
rect 8677 5525 8686 5655
rect 8612 5516 8686 5525
rect 10270 5655 10344 5664
rect 10270 5525 10279 5655
rect 10335 5525 10344 5655
rect 10270 5516 10344 5525
rect 11468 5456 11524 7380
rect 11676 7331 11732 7380
rect 12906 7369 12980 7378
rect 11662 7322 11736 7331
rect 11662 7192 11671 7322
rect 11727 7192 11736 7322
rect 12906 7239 12915 7369
rect 12971 7239 12980 7369
rect 15043 7341 15049 7457
rect 15101 7424 15139 7457
rect 15267 7470 15323 7834
rect 15482 7652 15536 8128
rect 15455 7646 15583 7652
rect 15455 7594 15461 7646
rect 15577 7594 15583 7646
rect 15455 7588 15583 7594
rect 15267 7464 15369 7470
rect 15267 7428 15311 7464
rect 15101 7341 15107 7424
rect 15305 7348 15311 7428
rect 15363 7348 15369 7464
rect 15305 7342 15369 7348
rect 15043 7335 15107 7341
rect 12906 7230 12980 7239
rect 11662 7183 11736 7192
rect 11573 6790 11647 6799
rect 11573 6734 11582 6790
rect 11638 6734 11647 6790
rect 11573 6725 11647 6734
rect 11576 6535 11635 6725
rect 11571 6529 11635 6535
rect 11571 6477 11577 6529
rect 11629 6477 11635 6529
rect 11571 6471 11635 6477
rect 11465 5447 11539 5456
rect 11465 5317 11474 5447
rect 11530 5317 11539 5447
rect 11465 5308 11539 5317
rect 8478 4499 8552 4508
rect 8478 4369 8487 4499
rect 8543 4369 8552 4499
rect 8478 4360 8552 4369
rect 8612 4499 8686 4508
rect 8612 4369 8621 4499
rect 8677 4369 8686 4499
rect 8612 4360 8686 4369
rect 10270 4499 10344 4508
rect 10270 4369 10279 4499
rect 10335 4369 10344 4499
rect 10270 4360 10344 4369
rect 8478 3343 8552 3352
rect 8478 3213 8487 3343
rect 8543 3213 8552 3343
rect 8478 3204 8552 3213
rect 8612 3343 8686 3352
rect 8612 3213 8621 3343
rect 8677 3213 8686 3343
rect 8612 3204 8686 3213
rect 10270 3343 10344 3352
rect 10270 3213 10279 3343
rect 10335 3213 10344 3343
rect 10270 3204 10344 3213
rect 11676 3004 11732 7183
rect 13812 7169 13886 7178
rect 13812 7039 13821 7169
rect 13877 7039 13886 7169
rect 13812 7030 13886 7039
rect 12146 6855 12220 6864
rect 12146 6725 12155 6855
rect 12211 6725 12220 6855
rect 12146 6716 12220 6725
rect 12314 6855 12388 6864
rect 12314 6725 12323 6855
rect 12379 6725 12388 6855
rect 12314 6716 12388 6725
rect 12447 6855 12521 6864
rect 12447 6725 12456 6855
rect 12512 6725 12521 6855
rect 12447 6716 12521 6725
rect 13363 6855 13437 6864
rect 13363 6725 13372 6855
rect 13428 6725 13437 6855
rect 13363 6716 13437 6725
rect 14279 6855 14353 6864
rect 14279 6725 14288 6855
rect 14344 6725 14353 6855
rect 14279 6716 14353 6725
rect 14413 6855 14487 6864
rect 14413 6725 14422 6855
rect 14478 6725 14487 6855
rect 14413 6716 14487 6725
rect 14654 6855 14728 6864
rect 14654 6725 14663 6855
rect 14719 6725 14728 6855
rect 14654 6716 14728 6725
rect 14788 6855 14862 6864
rect 14788 6725 14797 6855
rect 14853 6725 14862 6855
rect 14788 6716 14862 6725
rect 15562 6855 15636 6864
rect 15562 6725 15571 6855
rect 15627 6725 15636 6855
rect 15562 6716 15636 6725
rect 15696 6855 15770 6864
rect 15696 6725 15705 6855
rect 15761 6725 15770 6855
rect 15696 6716 15770 6725
rect 12501 5845 12629 5851
rect 12501 5793 12507 5845
rect 12623 5793 12629 5845
rect 12501 5787 12629 5793
rect 11894 5418 12042 5427
rect 11894 5362 11903 5418
rect 12033 5362 12042 5418
rect 11894 5353 11939 5362
rect 11933 5287 11939 5353
rect 11991 5353 12042 5362
rect 11991 5287 11997 5353
rect 11933 4247 11997 5287
rect 12536 4695 12594 5787
rect 13586 5655 13660 5664
rect 13586 5525 13595 5655
rect 13651 5525 13660 5655
rect 13586 5516 13660 5525
rect 15244 5655 15318 5664
rect 15244 5525 15253 5655
rect 15309 5525 15318 5655
rect 15244 5516 15318 5525
rect 15378 5655 15452 5664
rect 15378 5525 15387 5655
rect 15443 5525 15452 5655
rect 15378 5516 15452 5525
rect 12501 4689 12629 4695
rect 12501 4637 12507 4689
rect 12623 4637 12629 4689
rect 12501 4631 12629 4637
rect 11933 4131 11939 4247
rect 11991 4131 11997 4247
rect 11674 2998 11738 3004
rect 11674 2882 11680 2998
rect 11732 2882 11738 2998
rect 11674 2876 11738 2882
rect 8478 2187 8552 2196
rect 8478 2057 8487 2187
rect 8543 2057 8552 2187
rect 8478 2048 8552 2057
rect 8612 2187 8686 2196
rect 8612 2057 8621 2187
rect 8677 2057 8686 2187
rect 8612 2048 8686 2057
rect 10270 2187 10344 2196
rect 10270 2057 10279 2187
rect 10335 2057 10344 2187
rect 10270 2048 10344 2057
rect 11933 1935 11997 4131
rect 12536 3539 12594 4631
rect 13586 4499 13660 4508
rect 13586 4369 13595 4499
rect 13651 4369 13660 4499
rect 13586 4360 13660 4369
rect 15244 4499 15318 4508
rect 15244 4369 15253 4499
rect 15309 4369 15318 4499
rect 15244 4360 15318 4369
rect 15378 4499 15452 4508
rect 15378 4369 15387 4499
rect 15443 4369 15452 4499
rect 15378 4360 15452 4369
rect 12501 3533 12629 3539
rect 12501 3481 12507 3533
rect 12623 3481 12629 3533
rect 12501 3475 12629 3481
rect 12536 2383 12594 3475
rect 13586 3343 13660 3352
rect 13586 3213 13595 3343
rect 13651 3213 13660 3343
rect 13586 3204 13660 3213
rect 15244 3343 15318 3352
rect 15244 3213 15253 3343
rect 15309 3213 15318 3343
rect 15244 3204 15318 3213
rect 15378 3343 15452 3352
rect 15378 3213 15387 3343
rect 15443 3213 15452 3343
rect 15378 3204 15452 3213
rect 12501 2377 12629 2383
rect 12501 2325 12507 2377
rect 12623 2325 12629 2377
rect 12501 2319 12629 2325
rect 11933 1819 11939 1935
rect 11991 1819 11997 1935
rect 8478 1031 8552 1040
rect 8478 901 8487 1031
rect 8543 901 8552 1031
rect 8478 892 8552 901
rect 8612 1031 8686 1040
rect 8612 901 8621 1031
rect 8677 901 8686 1031
rect 8612 892 8686 901
rect 10270 1031 10344 1040
rect 10270 901 10279 1031
rect 10335 901 10344 1031
rect 10270 892 10344 901
rect 11933 779 11997 1819
rect 12536 1227 12594 2319
rect 13586 2187 13660 2196
rect 13586 2057 13595 2187
rect 13651 2057 13660 2187
rect 13586 2048 13660 2057
rect 15244 2187 15318 2196
rect 15244 2057 15253 2187
rect 15309 2057 15318 2187
rect 15244 2048 15318 2057
rect 15378 2187 15452 2196
rect 15378 2057 15387 2187
rect 15443 2057 15452 2187
rect 15378 2048 15452 2057
rect 12501 1221 12629 1227
rect 12501 1169 12507 1221
rect 12623 1169 12629 1221
rect 12501 1163 12629 1169
rect 13586 1031 13660 1040
rect 13586 901 13595 1031
rect 13651 901 13660 1031
rect 13586 892 13660 901
rect 15244 1031 15318 1040
rect 15244 901 15253 1031
rect 15309 901 15318 1031
rect 15244 892 15318 901
rect 15378 1031 15452 1040
rect 15378 901 15387 1031
rect 15443 901 15452 1031
rect 15378 892 15452 901
rect 11933 663 11939 779
rect 11991 663 11997 779
rect 11933 657 11997 663
rect 8100 -646 8106 -408
rect 8396 -646 8402 -408
rect 8100 -652 8402 -646
<< via2 >>
rect 3649 11307 3779 11309
rect 3649 11255 3651 11307
rect 3651 11255 3777 11307
rect 3777 11255 3779 11307
rect 3649 11253 3779 11255
rect 4721 11307 4851 11309
rect 4721 11255 4723 11307
rect 4723 11255 4849 11307
rect 4849 11255 4851 11307
rect 4721 11253 4851 11255
rect 8083 11192 8139 11194
rect 8083 11066 8085 11192
rect 8085 11066 8137 11192
rect 8137 11066 8139 11192
rect 8083 11064 8139 11066
rect 9799 11192 9855 11194
rect 9799 11066 9801 11192
rect 9801 11066 9853 11192
rect 9853 11066 9855 11192
rect 9799 11064 9855 11066
rect 1082 10711 1138 10713
rect 1082 10585 1084 10711
rect 1084 10585 1136 10711
rect 1136 10585 1138 10711
rect 1082 10583 1138 10585
rect 1218 10711 1274 10713
rect 1218 10585 1220 10711
rect 1220 10585 1272 10711
rect 1272 10585 1274 10711
rect 1218 10583 1274 10585
rect 2076 10711 2132 10713
rect 2076 10585 2078 10711
rect 2078 10585 2130 10711
rect 2130 10585 2132 10711
rect 2076 10583 2132 10585
rect 3792 10711 3848 10713
rect 3792 10585 3794 10711
rect 3794 10585 3846 10711
rect 3846 10585 3848 10711
rect 3792 10583 3848 10585
rect 4650 10711 4706 10713
rect 4650 10585 4652 10711
rect 4652 10585 4704 10711
rect 4704 10585 4706 10711
rect 4650 10583 4706 10585
rect 6366 10711 6422 10713
rect 6366 10585 6368 10711
rect 6368 10585 6420 10711
rect 6420 10585 6422 10711
rect 6366 10583 6422 10585
rect 7225 10711 7281 10713
rect 7225 10585 7227 10711
rect 7227 10585 7279 10711
rect 7279 10585 7281 10711
rect 7225 10583 7281 10585
rect 8113 10589 8382 10709
rect 3649 10151 3779 10153
rect 3649 10099 3651 10151
rect 3651 10099 3777 10151
rect 3777 10099 3779 10151
rect 3649 10097 3779 10099
rect 4721 10151 4851 10153
rect 4721 10099 4723 10151
rect 4723 10099 4849 10151
rect 4849 10099 4851 10151
rect 4721 10097 4851 10099
rect 3649 9647 3779 9649
rect 3649 9595 3651 9647
rect 3651 9595 3777 9647
rect 3777 9595 3779 9647
rect 3649 9593 3779 9595
rect 4721 9647 4851 9649
rect 4721 9595 4723 9647
rect 4723 9595 4849 9647
rect 4849 9595 4851 9647
rect 4721 9593 4851 9595
rect 150 9083 206 9213
rect 1082 9211 1138 9213
rect 1082 9085 1084 9211
rect 1084 9085 1136 9211
rect 1136 9085 1138 9211
rect 1082 9083 1138 9085
rect 1218 9211 1274 9213
rect 1218 9085 1220 9211
rect 1220 9085 1272 9211
rect 1272 9085 1274 9211
rect 1218 9083 1274 9085
rect 4225 9137 4281 9139
rect 4225 9085 4227 9137
rect 4227 9085 4279 9137
rect 4279 9085 4281 9137
rect 4225 9083 4281 9085
rect 2077 8760 2133 8762
rect 2077 8634 2079 8760
rect 2079 8634 2131 8760
rect 2131 8634 2133 8760
rect 2077 8632 2133 8634
rect 3793 8760 3849 8762
rect 3793 8634 3795 8760
rect 3795 8634 3847 8760
rect 3847 8634 3849 8760
rect 3793 8632 3849 8634
rect 4651 8760 4707 8762
rect 4651 8634 4653 8760
rect 4653 8634 4705 8760
rect 4705 8634 4707 8760
rect 4651 8632 4707 8634
rect 3649 8497 3779 8499
rect 3649 8445 3651 8497
rect 3651 8445 3777 8497
rect 3777 8445 3779 8497
rect 3649 8443 3779 8445
rect 4721 8497 4851 8499
rect 4721 8445 4723 8497
rect 4723 8445 4849 8497
rect 4849 8445 4851 8497
rect 4721 8443 4851 8445
rect 7225 9211 7281 9213
rect 7225 9085 7227 9211
rect 7227 9085 7279 9211
rect 7279 9085 7281 9211
rect 7225 9083 7281 9085
rect 7359 9211 7415 9213
rect 7359 9085 7361 9211
rect 7361 9085 7413 9211
rect 7413 9085 7415 9211
rect 7359 9083 7415 9085
rect 7754 9083 7810 9213
rect 6367 8760 6423 8762
rect 6367 8634 6369 8760
rect 6369 8634 6421 8760
rect 6421 8634 6423 8760
rect 6367 8632 6423 8634
rect 7439 8609 7495 8739
rect 6943 8391 6999 8521
rect 5507 7926 5563 8056
rect 6951 7018 7007 7148
rect 7982 6725 8038 6855
rect 7982 5525 8038 5655
rect 7982 4369 8038 4499
rect 7982 3213 8038 3343
rect 7982 2057 8038 2187
rect 7982 901 8038 1031
rect 8941 10711 8997 10713
rect 8941 10585 8943 10711
rect 8943 10585 8995 10711
rect 8995 10585 8997 10711
rect 8941 10583 8997 10585
rect 10657 10711 10713 10713
rect 10657 10585 10659 10711
rect 10659 10585 10711 10711
rect 10711 10585 10713 10711
rect 10657 10583 10713 10585
rect 12373 10711 12429 10713
rect 12373 10585 12375 10711
rect 12375 10585 12427 10711
rect 12427 10585 12429 10711
rect 12373 10583 12429 10585
rect 13231 10711 13287 10713
rect 13231 10585 13233 10711
rect 13233 10585 13285 10711
rect 13285 10585 13287 10711
rect 13231 10583 13287 10585
rect 13364 10711 13420 10713
rect 13364 10585 13366 10711
rect 13366 10585 13418 10711
rect 13418 10585 13420 10711
rect 13364 10583 13420 10585
rect 10610 9491 10740 9547
rect 10462 9327 10518 9329
rect 10462 9275 10464 9327
rect 10464 9275 10516 9327
rect 10516 9275 10518 9327
rect 10462 9273 10518 9275
rect 10285 8868 10341 8998
rect 8337 8548 8393 8678
rect 10235 8676 10291 8678
rect 10235 8550 10237 8676
rect 10237 8550 10289 8676
rect 10289 8550 10291 8676
rect 10235 8548 10291 8550
rect 10355 8364 10411 8366
rect 10355 8238 10357 8364
rect 10357 8238 10409 8364
rect 10409 8238 10411 8364
rect 10355 8236 10411 8238
rect 8993 7171 9049 7173
rect 8993 7045 8995 7171
rect 8995 7045 9047 7171
rect 9047 7045 9049 7171
rect 8993 7043 9049 7045
rect 8861 6853 8917 6855
rect 8861 6727 8863 6853
rect 8863 6727 8915 6853
rect 8915 6727 8917 6853
rect 8861 6725 8917 6727
rect 10725 8707 10781 8709
rect 10725 8655 10727 8707
rect 10727 8655 10779 8707
rect 10779 8655 10781 8707
rect 10725 8653 10781 8655
rect 10941 9140 10997 9142
rect 10941 9014 10943 9140
rect 10943 9014 10995 9140
rect 10995 9014 10997 9140
rect 10941 9012 10997 9014
rect 11046 8918 11102 8920
rect 11046 8792 11048 8918
rect 11048 8792 11100 8918
rect 11100 8792 11102 8918
rect 11046 8790 11102 8792
rect 12304 9487 12434 9543
rect 13902 9489 14032 9545
rect 15411 9489 15541 9545
rect 11426 8890 11482 9020
rect 10814 8549 10870 8605
rect 11170 8549 11226 8605
rect 11880 9318 11936 9320
rect 11880 9266 11882 9318
rect 11882 9266 11934 9318
rect 11934 9266 11936 9318
rect 11880 9264 11936 9266
rect 11526 8549 11582 8605
rect 10625 8192 10681 8194
rect 10625 8140 10627 8192
rect 10627 8140 10679 8192
rect 10679 8140 10681 8192
rect 10625 8138 10681 8140
rect 10981 8192 11037 8194
rect 10981 8140 10983 8192
rect 10983 8140 11035 8192
rect 11035 8140 11037 8192
rect 10981 8138 11037 8140
rect 10896 7945 10952 8001
rect 11039 7988 11095 8044
rect 10346 7390 10402 7520
rect 11048 7846 11104 7902
rect 11348 8202 11404 8204
rect 11348 8150 11350 8202
rect 11350 8150 11402 8202
rect 11402 8150 11404 8202
rect 11348 8148 11404 8150
rect 11345 7848 11401 7904
rect 11402 7640 11458 7642
rect 11402 7588 11404 7640
rect 11404 7588 11456 7640
rect 11456 7588 11458 7640
rect 11402 7586 11458 7588
rect 13614 9179 13670 9181
rect 13614 9053 13616 9179
rect 13616 9053 13668 9179
rect 13668 9053 13670 9179
rect 13614 9051 13670 9053
rect 12693 9010 12749 9012
rect 12693 8884 12695 9010
rect 12695 8884 12747 9010
rect 12747 8884 12749 9010
rect 12693 8882 12749 8884
rect 12103 8676 12159 8678
rect 12103 8550 12105 8676
rect 12105 8550 12157 8676
rect 12157 8550 12159 8676
rect 12103 8548 12159 8550
rect 12239 8676 12295 8678
rect 12239 8550 12241 8676
rect 12241 8550 12293 8676
rect 12293 8550 12295 8676
rect 12239 8548 12295 8550
rect 13155 8676 13211 8678
rect 13155 8550 13157 8676
rect 13157 8550 13209 8676
rect 13209 8550 13211 8676
rect 13155 8548 13211 8550
rect 11756 8166 11812 8168
rect 11756 8114 11758 8166
rect 11758 8114 11810 8166
rect 11810 8114 11812 8166
rect 11756 8112 11812 8114
rect 11788 7976 11844 8032
rect 11933 7977 11989 8033
rect 11760 7640 11816 7642
rect 11760 7588 11762 7640
rect 11762 7588 11814 7640
rect 11814 7588 11816 7640
rect 11760 7586 11816 7588
rect 11917 7655 11973 7657
rect 11917 7603 11919 7655
rect 11919 7603 11971 7655
rect 11971 7603 11973 7655
rect 11917 7601 11973 7603
rect 12982 7980 13112 8036
rect 12561 7846 12617 7902
rect 13707 7850 13763 7906
rect 13461 7671 13517 7727
rect 14532 8894 14588 8896
rect 14532 8768 14534 8894
rect 14534 8768 14586 8894
rect 14586 8768 14588 8894
rect 14532 8766 14588 8768
rect 14071 8676 14127 8678
rect 14071 8550 14073 8676
rect 14073 8550 14125 8676
rect 14125 8550 14127 8676
rect 14071 8548 14127 8550
rect 14663 8676 14719 8678
rect 14663 8550 14665 8676
rect 14665 8550 14717 8676
rect 14717 8550 14719 8676
rect 14663 8548 14719 8550
rect 14797 8676 14853 8678
rect 14797 8550 14799 8676
rect 14799 8550 14851 8676
rect 14851 8550 14853 8676
rect 14797 8548 14853 8550
rect 14176 7676 14232 7732
rect 15081 7973 15137 8029
rect 15571 8676 15627 8678
rect 15571 8550 15573 8676
rect 15573 8550 15625 8676
rect 15625 8550 15627 8676
rect 15571 8548 15627 8550
rect 15703 8676 15759 8678
rect 15703 8550 15705 8676
rect 15705 8550 15757 8676
rect 15757 8550 15759 8676
rect 15703 8548 15759 8550
rect 15266 7843 15322 7899
rect 9175 7335 9231 7337
rect 9175 7209 9177 7335
rect 9177 7209 9229 7335
rect 9229 7209 9231 7335
rect 9175 7207 9231 7209
rect 9529 7335 9585 7337
rect 9529 7209 9531 7335
rect 9531 7209 9583 7335
rect 9583 7209 9585 7335
rect 9529 7207 9585 7209
rect 9885 7335 9941 7337
rect 9885 7209 9887 7335
rect 9887 7209 9939 7335
rect 9939 7209 9941 7335
rect 9885 7207 9941 7209
rect 10241 7335 10297 7337
rect 10241 7209 10243 7335
rect 10243 7209 10295 7335
rect 10295 7209 10297 7335
rect 10241 7207 10297 7209
rect 10597 7335 10653 7337
rect 10597 7209 10599 7335
rect 10599 7209 10651 7335
rect 10651 7209 10653 7335
rect 10597 7207 10653 7209
rect 9351 7171 9407 7173
rect 9351 7045 9353 7171
rect 9353 7045 9405 7171
rect 9405 7045 9407 7171
rect 9351 7043 9407 7045
rect 9707 7171 9763 7173
rect 9707 7045 9709 7171
rect 9709 7045 9761 7171
rect 9761 7045 9763 7171
rect 9707 7043 9763 7045
rect 10063 7171 10119 7173
rect 10063 7045 10065 7171
rect 10065 7045 10117 7171
rect 10117 7045 10119 7171
rect 10063 7043 10119 7045
rect 10419 7171 10475 7173
rect 10419 7045 10421 7171
rect 10421 7045 10473 7171
rect 10473 7045 10475 7171
rect 10419 7043 10475 7045
rect 10775 7171 10831 7173
rect 10775 7045 10777 7171
rect 10777 7045 10829 7171
rect 10829 7045 10831 7171
rect 10775 7043 10831 7045
rect 10860 6737 10916 6793
rect 11216 6738 11272 6794
rect 8487 5653 8543 5655
rect 8487 5527 8489 5653
rect 8489 5527 8541 5653
rect 8541 5527 8543 5653
rect 8487 5525 8543 5527
rect 8621 5653 8677 5655
rect 8621 5527 8623 5653
rect 8623 5527 8675 5653
rect 8675 5527 8677 5653
rect 8621 5525 8677 5527
rect 10279 5653 10335 5655
rect 10279 5527 10281 5653
rect 10281 5527 10333 5653
rect 10333 5527 10335 5653
rect 10279 5525 10335 5527
rect 11671 7192 11727 7322
rect 12915 7367 12971 7369
rect 12915 7241 12917 7367
rect 12917 7241 12969 7367
rect 12969 7241 12971 7367
rect 12915 7239 12971 7241
rect 11582 6734 11638 6790
rect 11474 5317 11530 5447
rect 8487 4497 8543 4499
rect 8487 4371 8489 4497
rect 8489 4371 8541 4497
rect 8541 4371 8543 4497
rect 8487 4369 8543 4371
rect 8621 4497 8677 4499
rect 8621 4371 8623 4497
rect 8623 4371 8675 4497
rect 8675 4371 8677 4497
rect 8621 4369 8677 4371
rect 10279 4497 10335 4499
rect 10279 4371 10281 4497
rect 10281 4371 10333 4497
rect 10333 4371 10335 4497
rect 10279 4369 10335 4371
rect 8487 3341 8543 3343
rect 8487 3215 8489 3341
rect 8489 3215 8541 3341
rect 8541 3215 8543 3341
rect 8487 3213 8543 3215
rect 8621 3341 8677 3343
rect 8621 3215 8623 3341
rect 8623 3215 8675 3341
rect 8675 3215 8677 3341
rect 8621 3213 8677 3215
rect 10279 3341 10335 3343
rect 10279 3215 10281 3341
rect 10281 3215 10333 3341
rect 10333 3215 10335 3341
rect 10279 3213 10335 3215
rect 13821 7167 13877 7169
rect 13821 7041 13823 7167
rect 13823 7041 13875 7167
rect 13875 7041 13877 7167
rect 13821 7039 13877 7041
rect 12155 6853 12211 6855
rect 12155 6727 12157 6853
rect 12157 6727 12209 6853
rect 12209 6727 12211 6853
rect 12155 6725 12211 6727
rect 12323 6853 12379 6855
rect 12323 6727 12325 6853
rect 12325 6727 12377 6853
rect 12377 6727 12379 6853
rect 12323 6725 12379 6727
rect 12456 6853 12512 6855
rect 12456 6727 12458 6853
rect 12458 6727 12510 6853
rect 12510 6727 12512 6853
rect 12456 6725 12512 6727
rect 13372 6853 13428 6855
rect 13372 6727 13374 6853
rect 13374 6727 13426 6853
rect 13426 6727 13428 6853
rect 13372 6725 13428 6727
rect 14288 6853 14344 6855
rect 14288 6727 14290 6853
rect 14290 6727 14342 6853
rect 14342 6727 14344 6853
rect 14288 6725 14344 6727
rect 14422 6853 14478 6855
rect 14422 6727 14424 6853
rect 14424 6727 14476 6853
rect 14476 6727 14478 6853
rect 14422 6725 14478 6727
rect 14663 6853 14719 6855
rect 14663 6727 14665 6853
rect 14665 6727 14717 6853
rect 14717 6727 14719 6853
rect 14663 6725 14719 6727
rect 14797 6853 14853 6855
rect 14797 6727 14799 6853
rect 14799 6727 14851 6853
rect 14851 6727 14853 6853
rect 14797 6725 14853 6727
rect 15571 6853 15627 6855
rect 15571 6727 15573 6853
rect 15573 6727 15625 6853
rect 15625 6727 15627 6853
rect 15571 6725 15627 6727
rect 15705 6853 15761 6855
rect 15705 6727 15707 6853
rect 15707 6727 15759 6853
rect 15759 6727 15761 6853
rect 15705 6725 15761 6727
rect 11903 5416 12033 5418
rect 11903 5364 11905 5416
rect 11905 5364 12031 5416
rect 12031 5364 12033 5416
rect 11903 5362 11939 5364
rect 11939 5362 11991 5364
rect 11991 5362 12033 5364
rect 13595 5653 13651 5655
rect 13595 5527 13597 5653
rect 13597 5527 13649 5653
rect 13649 5527 13651 5653
rect 13595 5525 13651 5527
rect 15253 5653 15309 5655
rect 15253 5527 15255 5653
rect 15255 5527 15307 5653
rect 15307 5527 15309 5653
rect 15253 5525 15309 5527
rect 15387 5653 15443 5655
rect 15387 5527 15389 5653
rect 15389 5527 15441 5653
rect 15441 5527 15443 5653
rect 15387 5525 15443 5527
rect 8487 2185 8543 2187
rect 8487 2059 8489 2185
rect 8489 2059 8541 2185
rect 8541 2059 8543 2185
rect 8487 2057 8543 2059
rect 8621 2185 8677 2187
rect 8621 2059 8623 2185
rect 8623 2059 8675 2185
rect 8675 2059 8677 2185
rect 8621 2057 8677 2059
rect 10279 2185 10335 2187
rect 10279 2059 10281 2185
rect 10281 2059 10333 2185
rect 10333 2059 10335 2185
rect 10279 2057 10335 2059
rect 13595 4497 13651 4499
rect 13595 4371 13597 4497
rect 13597 4371 13649 4497
rect 13649 4371 13651 4497
rect 13595 4369 13651 4371
rect 15253 4497 15309 4499
rect 15253 4371 15255 4497
rect 15255 4371 15307 4497
rect 15307 4371 15309 4497
rect 15253 4369 15309 4371
rect 15387 4497 15443 4499
rect 15387 4371 15389 4497
rect 15389 4371 15441 4497
rect 15441 4371 15443 4497
rect 15387 4369 15443 4371
rect 13595 3341 13651 3343
rect 13595 3215 13597 3341
rect 13597 3215 13649 3341
rect 13649 3215 13651 3341
rect 13595 3213 13651 3215
rect 15253 3341 15309 3343
rect 15253 3215 15255 3341
rect 15255 3215 15307 3341
rect 15307 3215 15309 3341
rect 15253 3213 15309 3215
rect 15387 3341 15443 3343
rect 15387 3215 15389 3341
rect 15389 3215 15441 3341
rect 15441 3215 15443 3341
rect 15387 3213 15443 3215
rect 8487 1029 8543 1031
rect 8487 903 8489 1029
rect 8489 903 8541 1029
rect 8541 903 8543 1029
rect 8487 901 8543 903
rect 8621 1029 8677 1031
rect 8621 903 8623 1029
rect 8623 903 8675 1029
rect 8675 903 8677 1029
rect 8621 901 8677 903
rect 10279 1029 10335 1031
rect 10279 903 10281 1029
rect 10281 903 10333 1029
rect 10333 903 10335 1029
rect 10279 901 10335 903
rect 13595 2185 13651 2187
rect 13595 2059 13597 2185
rect 13597 2059 13649 2185
rect 13649 2059 13651 2185
rect 13595 2057 13651 2059
rect 15253 2185 15309 2187
rect 15253 2059 15255 2185
rect 15255 2059 15307 2185
rect 15307 2059 15309 2185
rect 15253 2057 15309 2059
rect 15387 2185 15443 2187
rect 15387 2059 15389 2185
rect 15389 2059 15441 2185
rect 15441 2059 15443 2185
rect 15387 2057 15443 2059
rect 13595 1029 13651 1031
rect 13595 903 13597 1029
rect 13597 903 13649 1029
rect 13649 903 13651 1029
rect 13595 901 13651 903
rect 15253 1029 15309 1031
rect 15253 903 15255 1029
rect 15255 903 15307 1029
rect 15307 903 15309 1029
rect 15253 901 15309 903
rect 15387 1029 15443 1031
rect 15387 903 15389 1029
rect 15389 903 15441 1029
rect 15441 903 15443 1029
rect 15387 901 15443 903
<< metal3 >>
rect 3640 11311 3788 11318
rect 4712 11311 4860 11318
rect 3640 11309 4860 11311
rect 3640 11253 3649 11309
rect 3779 11253 4721 11309
rect 4851 11253 4860 11309
rect 3640 11251 4860 11253
rect 3640 11244 3788 11251
rect 4712 11244 4860 11251
rect 8074 11194 8148 11203
rect 8074 11064 8083 11194
rect 8139 11064 8148 11194
rect 8074 11055 8148 11064
rect 9790 11194 9864 11203
rect 9790 11064 9799 11194
rect 9855 11064 9864 11194
rect 9790 11055 9864 11064
rect 1073 10713 13429 10722
rect 1073 10583 1082 10713
rect 1138 10583 1218 10713
rect 1274 10583 2076 10713
rect 2132 10583 3792 10713
rect 3848 10583 4650 10713
rect 4706 10583 6366 10713
rect 6422 10583 7225 10713
rect 7281 10709 8941 10713
rect 7281 10589 8113 10709
rect 8382 10589 8941 10709
rect 7281 10583 8941 10589
rect 8997 10583 10657 10713
rect 10713 10583 12373 10713
rect 12429 10583 13231 10713
rect 13287 10583 13364 10713
rect 13420 10583 13429 10713
rect 1073 10574 13429 10583
rect 3640 10155 3788 10162
rect 4712 10155 4860 10162
rect 3640 10153 4860 10155
rect 3640 10097 3649 10153
rect 3779 10097 4721 10153
rect 4851 10097 4860 10153
rect 3640 10095 4860 10097
rect 3640 10088 3788 10095
rect 4712 10088 4860 10095
rect 3640 9651 3788 9658
rect 4712 9651 4860 9658
rect 3640 9649 4860 9651
rect 3640 9593 3649 9649
rect 3779 9593 4721 9649
rect 4851 9593 4860 9649
rect 3640 9591 4860 9593
rect 3640 9584 3788 9591
rect 4712 9584 4860 9591
rect 10601 9548 10749 9556
rect 12295 9548 12443 9552
rect 13893 9549 14041 9554
rect 15402 9549 15550 9554
rect 13893 9548 15550 9549
rect 10601 9547 15550 9548
rect 10601 9491 10610 9547
rect 10740 9545 15550 9547
rect 10740 9543 13902 9545
rect 10740 9491 12304 9543
rect 10601 9488 12304 9491
rect 10601 9482 10749 9488
rect 12295 9487 12304 9488
rect 12434 9489 13902 9543
rect 14032 9489 15411 9545
rect 15541 9489 15550 9545
rect 12434 9488 14041 9489
rect 12434 9487 12443 9488
rect 12295 9478 12443 9487
rect 13893 9480 14041 9488
rect 15402 9480 15550 9489
rect 10453 9329 10527 9338
rect 10453 9273 10462 9329
rect 10518 9327 10527 9329
rect 11871 9327 11945 9329
rect 10518 9320 11945 9327
rect 10518 9273 11880 9320
rect 10453 9264 11880 9273
rect 11936 9264 11945 9320
rect 10513 9261 11945 9264
rect 11871 9255 11945 9261
rect 141 9213 7819 9222
rect 141 9083 150 9213
rect 206 9083 1082 9213
rect 1138 9083 1218 9213
rect 1274 9139 7225 9213
rect 1274 9083 4225 9139
rect 4281 9083 7225 9139
rect 7281 9083 7359 9213
rect 7415 9083 7754 9213
rect 7810 9083 7819 9213
rect 13605 9181 13679 9190
rect 13605 9155 13614 9181
rect 10982 9151 13614 9155
rect 141 9074 7819 9083
rect 10932 9142 13614 9151
rect 10932 9012 10941 9142
rect 10997 9095 13614 9142
rect 10997 9012 11006 9095
rect 13605 9051 13614 9095
rect 13670 9051 13679 9181
rect 13605 9042 13679 9051
rect 10276 8998 10350 9007
rect 10932 9003 11006 9012
rect 11417 9020 11491 9029
rect 10276 8868 10285 8998
rect 10341 8927 10350 8998
rect 11037 8927 11111 8929
rect 10341 8920 11111 8927
rect 10341 8868 11046 8920
rect 10276 8867 11046 8868
rect 10276 8859 10350 8867
rect 11037 8790 11046 8867
rect 11102 8813 11111 8920
rect 11417 8890 11426 9020
rect 11482 8995 11491 9020
rect 12684 9012 12758 9021
rect 12684 8995 12693 9012
rect 11482 8935 12693 8995
rect 11482 8890 11491 8935
rect 11417 8881 11491 8890
rect 12684 8882 12693 8935
rect 12749 8882 12758 9012
rect 12684 8873 12758 8882
rect 14523 8896 14597 8905
rect 14523 8813 14532 8896
rect 11102 8790 14532 8813
rect 11037 8781 14532 8790
rect 2068 8762 2142 8771
rect 2068 8632 2077 8762
rect 2133 8683 2142 8762
rect 3784 8762 3858 8771
rect 3784 8683 3793 8762
rect 2133 8632 3793 8683
rect 3849 8632 3858 8762
rect 2068 8623 3858 8632
rect 4642 8762 4716 8771
rect 4642 8632 4651 8762
rect 4707 8683 4716 8762
rect 6358 8762 6432 8771
rect 6358 8683 6367 8762
rect 4707 8632 6367 8683
rect 6423 8683 6432 8762
rect 11038 8766 14532 8781
rect 14588 8766 14597 8896
rect 11038 8757 14597 8766
rect 11038 8753 14583 8757
rect 7430 8739 7504 8748
rect 7430 8683 7439 8739
rect 6423 8632 7439 8683
rect 4642 8623 7439 8632
rect 7430 8609 7439 8623
rect 7495 8609 7504 8739
rect 10716 8709 10790 8718
rect 10716 8687 10725 8709
rect 7430 8600 7504 8609
rect 8328 8678 10725 8687
rect 8328 8548 8337 8678
rect 8393 8548 10235 8678
rect 10291 8653 10725 8678
rect 10781 8687 10790 8709
rect 10781 8678 15768 8687
rect 10781 8653 12103 8678
rect 10291 8605 12103 8653
rect 10291 8549 10814 8605
rect 10870 8549 11170 8605
rect 11226 8549 11526 8605
rect 11582 8549 12103 8605
rect 10291 8548 12103 8549
rect 12159 8548 12239 8678
rect 12295 8548 13155 8678
rect 13211 8548 14071 8678
rect 14127 8548 14663 8678
rect 14719 8548 14797 8678
rect 14853 8548 15571 8678
rect 15627 8548 15703 8678
rect 15759 8548 15768 8678
rect 8328 8539 15768 8548
rect 6934 8521 7008 8530
rect 3640 8501 3788 8508
rect 4712 8501 4860 8508
rect 6934 8501 6943 8521
rect 3640 8499 6943 8501
rect 3640 8443 3649 8499
rect 3779 8443 4721 8499
rect 4851 8443 6943 8499
rect 3640 8441 6943 8443
rect 3640 8434 3788 8441
rect 4712 8434 4860 8441
rect 6934 8391 6943 8441
rect 6999 8391 7008 8521
rect 6934 8382 7008 8391
rect 10346 8366 10420 8375
rect 10346 8236 10355 8366
rect 10411 8236 10420 8366
rect 10346 8227 10420 8236
rect 11339 8204 11807 8213
rect 10616 8194 11046 8203
rect 10616 8138 10625 8194
rect 10681 8138 10981 8194
rect 11037 8138 11046 8194
rect 11339 8148 11348 8204
rect 11404 8177 11807 8204
rect 11404 8168 11821 8177
rect 11404 8148 11756 8168
rect 11339 8139 11756 8148
rect 10616 8129 11046 8138
rect 11747 8112 11756 8139
rect 11812 8112 11821 8168
rect 11747 8103 11821 8112
rect 5498 8056 5572 8065
rect 5498 7926 5507 8056
rect 5563 8008 5572 8056
rect 11030 8044 11104 8053
rect 10887 8008 10961 8010
rect 5563 8001 10961 8008
rect 5563 7945 10896 8001
rect 10952 7945 10961 8001
rect 11030 7988 11039 8044
rect 11095 8039 11104 8044
rect 11779 8039 11853 8041
rect 11095 8032 11853 8039
rect 11095 7988 11788 8032
rect 11030 7979 11788 7988
rect 11779 7976 11788 7979
rect 11844 7976 11853 8032
rect 11779 7967 11853 7976
rect 11924 8035 11998 8042
rect 12973 8036 13121 8045
rect 12973 8035 12982 8036
rect 11924 8033 12982 8035
rect 11924 7977 11933 8033
rect 11989 7980 12982 8033
rect 13112 8035 13121 8036
rect 15072 8035 15146 8038
rect 13112 8029 15146 8035
rect 13112 7980 15081 8029
rect 11989 7977 15081 7980
rect 11924 7975 15081 7977
rect 11924 7968 11998 7975
rect 12973 7971 13121 7975
rect 15072 7973 15081 7975
rect 15137 7973 15146 8029
rect 15072 7964 15146 7973
rect 5563 7937 10961 7945
rect 5563 7926 5572 7937
rect 10887 7936 10961 7937
rect 5498 7917 5572 7926
rect 11336 7911 11410 7913
rect 11039 7907 11410 7911
rect 12552 7907 12626 7911
rect 13698 7907 13772 7915
rect 11039 7906 13772 7907
rect 11039 7904 13707 7906
rect 11039 7902 11345 7904
rect 11039 7846 11048 7902
rect 11104 7848 11345 7902
rect 11401 7902 13707 7904
rect 11401 7848 12561 7902
rect 11104 7847 12561 7848
rect 11104 7846 11113 7847
rect 11039 7837 11113 7846
rect 11336 7839 11410 7847
rect 12552 7846 12561 7847
rect 12617 7850 13707 7902
rect 13763 7904 13772 7906
rect 15257 7904 15331 7908
rect 13763 7899 15331 7904
rect 13763 7850 15266 7899
rect 12617 7847 15266 7850
rect 12617 7846 12626 7847
rect 12552 7837 12626 7846
rect 13698 7844 15266 7847
rect 13698 7841 13772 7844
rect 15257 7843 15266 7844
rect 15322 7843 15331 7899
rect 15257 7834 15331 7843
rect 13452 7727 13526 7736
rect 13452 7721 13461 7727
rect 11909 7671 13461 7721
rect 13517 7721 13526 7727
rect 14167 7732 14241 7741
rect 14167 7721 14176 7732
rect 13517 7676 14176 7721
rect 14232 7676 14241 7732
rect 13517 7671 14241 7676
rect 11909 7667 14241 7671
rect 11909 7666 14202 7667
rect 11908 7661 14202 7666
rect 11908 7657 11982 7661
rect 11393 7642 11825 7651
rect 11393 7586 11402 7642
rect 11458 7586 11760 7642
rect 11816 7586 11825 7642
rect 11908 7601 11917 7657
rect 11973 7601 11982 7657
rect 11908 7592 11982 7601
rect 11393 7577 11825 7586
rect 10337 7520 10411 7529
rect 10337 7390 10346 7520
rect 10402 7390 10411 7520
rect 10337 7346 10411 7390
rect 12906 7369 12980 7378
rect 9166 7337 10662 7346
rect 9166 7207 9175 7337
rect 9231 7286 9529 7337
rect 9231 7207 9240 7286
rect 9166 7198 9240 7207
rect 9520 7207 9529 7286
rect 9585 7286 9885 7337
rect 9585 7207 9594 7286
rect 9520 7198 9594 7207
rect 9876 7207 9885 7286
rect 9941 7286 10241 7337
rect 9941 7207 9950 7286
rect 9876 7198 9950 7207
rect 10232 7207 10241 7286
rect 10297 7286 10597 7337
rect 10297 7207 10306 7286
rect 10232 7198 10306 7207
rect 10588 7207 10597 7286
rect 10653 7207 10662 7337
rect 10588 7198 10662 7207
rect 11662 7322 11736 7331
rect 11662 7192 11671 7322
rect 11727 7314 11736 7322
rect 12906 7314 12915 7369
rect 11727 7254 12915 7314
rect 11727 7192 11736 7254
rect 12906 7239 12915 7254
rect 12971 7239 12980 7369
rect 12906 7230 12980 7239
rect 11662 7183 11736 7192
rect 8984 7173 9058 7182
rect 6942 7148 7016 7157
rect 6942 7018 6951 7148
rect 7007 7094 7016 7148
rect 8984 7094 8993 7173
rect 7007 7043 8993 7094
rect 9049 7094 9058 7173
rect 9342 7173 9416 7182
rect 9342 7094 9351 7173
rect 9049 7043 9351 7094
rect 9407 7094 9416 7173
rect 9698 7173 9772 7182
rect 9698 7094 9707 7173
rect 9407 7043 9707 7094
rect 9763 7094 9772 7173
rect 10054 7173 10128 7182
rect 10054 7094 10063 7173
rect 9763 7043 10063 7094
rect 10119 7094 10128 7173
rect 10410 7173 10484 7182
rect 10410 7094 10419 7173
rect 10119 7043 10419 7094
rect 10475 7094 10484 7173
rect 10766 7173 10840 7182
rect 10766 7094 10775 7173
rect 10475 7043 10775 7094
rect 10831 7094 10840 7173
rect 13812 7169 13886 7178
rect 13812 7094 13821 7169
rect 10831 7043 13821 7094
rect 7007 7039 13821 7043
rect 13877 7039 13886 7169
rect 7007 7034 13886 7039
rect 7007 7018 7016 7034
rect 13812 7030 13886 7034
rect 6942 7009 7016 7018
rect 7973 6855 15770 6864
rect 7973 6725 7982 6855
rect 8038 6725 8861 6855
rect 8917 6794 12155 6855
rect 8917 6793 11216 6794
rect 8917 6737 10860 6793
rect 10916 6738 11216 6793
rect 11272 6790 12155 6794
rect 11272 6738 11582 6790
rect 10916 6737 11582 6738
rect 8917 6734 11582 6737
rect 11638 6734 12155 6790
rect 8917 6725 12155 6734
rect 12211 6725 12323 6855
rect 12379 6725 12456 6855
rect 12512 6725 13372 6855
rect 13428 6725 14288 6855
rect 14344 6725 14422 6855
rect 14478 6725 14663 6855
rect 14719 6725 14797 6855
rect 14853 6725 15571 6855
rect 15627 6725 15705 6855
rect 15761 6725 15770 6855
rect 7973 6716 15770 6725
rect 7973 5655 15452 5664
rect 7973 5525 7982 5655
rect 8038 5525 8487 5655
rect 8543 5525 8621 5655
rect 8677 5525 10279 5655
rect 10335 5525 13595 5655
rect 13651 5525 15253 5655
rect 15309 5525 15387 5655
rect 15443 5525 15452 5655
rect 7973 5516 15452 5525
rect 11465 5447 11539 5456
rect 11465 5317 11474 5447
rect 11530 5427 11539 5447
rect 11530 5418 12042 5427
rect 11530 5362 11903 5418
rect 12033 5362 12042 5418
rect 11530 5353 12042 5362
rect 11530 5317 11539 5353
rect 11465 5308 11539 5317
rect 7973 4499 15452 4508
rect 7973 4369 7982 4499
rect 8038 4369 8487 4499
rect 8543 4369 8621 4499
rect 8677 4369 10279 4499
rect 10335 4369 13595 4499
rect 13651 4369 15253 4499
rect 15309 4369 15387 4499
rect 15443 4369 15452 4499
rect 7973 4360 15452 4369
rect 7973 3343 15452 3352
rect 7973 3213 7982 3343
rect 8038 3213 8487 3343
rect 8543 3213 8621 3343
rect 8677 3213 10279 3343
rect 10335 3213 13595 3343
rect 13651 3213 15253 3343
rect 15309 3213 15387 3343
rect 15443 3213 15452 3343
rect 7973 3204 15452 3213
rect 7973 2187 15452 2196
rect 7973 2057 7982 2187
rect 8038 2057 8487 2187
rect 8543 2057 8621 2187
rect 8677 2057 10279 2187
rect 10335 2057 13595 2187
rect 13651 2057 15253 2187
rect 15309 2057 15387 2187
rect 15443 2057 15452 2187
rect 7973 2048 15452 2057
rect 7973 1031 15452 1040
rect 7973 901 7982 1031
rect 8038 901 8487 1031
rect 8543 901 8621 1031
rect 8677 901 10279 1031
rect 10335 901 13595 1031
rect 13651 901 15253 1031
rect 15309 901 15387 1031
rect 15443 901 15452 1031
rect 7973 892 15452 901
use sky130_fd_pr__nfet_g5v0d10v5_3DCHX4  sky130_fd_pr__nfet_g5v0d10v5_3DCHX4_0
timestamp 1712352531
transform 1 0 11965 0 1 2974
box -3515 -3039 3515 3039
use sky130_fd_pr__nfet_g5v0d10v5_62W3XE  sky130_fd_pr__nfet_g5v0d10v5_62W3XE_0
timestamp 1712352531
transform 1 0 15212 0 1 7049
box -586 -758 586 758
use sky130_fd_pr__nfet_g5v0d10v5_EC8RE7  sky130_fd_pr__nfet_g5v0d10v5_EC8RE7_1
timestamp 1712352531
transform 1 0 10536 0 1 7049
box -1712 -758 1712 758
use sky130_fd_pr__nfet_g5v0d10v5_QZVU2P  sky130_fd_pr__nfet_g5v0d10v5_QZVU2P_1
timestamp 1712352531
transform 1 0 4250 0 1 9046
box -3202 -758 3202 758
use sky130_fd_pr__nfet_g5v0d10v5_XZ4X25  sky130_fd_pr__nfet_g5v0d10v5_XZ4X25_0
timestamp 1712352531
transform 1 0 13400 0 1 7049
box -1115 -758 1115 758
use sky130_fd_pr__pfet_g5v0d10v5_7JLQGA  sky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0
timestamp 1712352531
transform 1 0 11198 0 1 8727
box -1030 -797 1030 797
use sky130_fd_pr__pfet_g5v0d10v5_75AJMX  sky130_fd_pr__pfet_g5v0d10v5_75AJMX_0
timestamp 1712352531
transform 1 0 7253 0 1 10703
box -6235 -797 6235 797
use sky130_fd_pr__pfet_g5v0d10v5_Y9J9EP  sky130_fd_pr__pfet_g5v0d10v5_Y9J9EP_0
timestamp 1712352531
transform 1 0 15212 0 1 8727
box -616 -797 616 797
use sky130_fd_pr__pfet_g5v0d10v5_Y9S9FP  sky130_fd_pr__pfet_g5v0d10v5_Y9S9FP_0
timestamp 1712352531
transform 1 0 13412 0 1 8727
box -1374 -797 1374 797
use sky130_fd_pr__res_xhigh_po_1p41_DVQADA  sky130_fd_pr__res_xhigh_po_1p41_DVQADA_0
timestamp 1712352531
transform 1 0 3845 0 1 4029
box -3898 -4082 3898 4082
<< labels >>
flabel metal2 123 7939 123 7939 0 FreeSans 1200 0 0 0 avss
port 8 nsew
flabel metal3 4681 9651 4681 9651 0 FreeSans 800 0 0 0 vn0
flabel metal3 7414 8683 7414 8683 0 FreeSans 800 0 0 0 vr
flabel comment s 1668 9043 1668 9043 0 FreeSans 800 0 0 0 dum
flabel comment s 2526 9043 2526 9043 0 FreeSans 800 0 0 0 Mn0
flabel comment s 3384 9043 3384 9043 0 FreeSans 800 0 0 0 Mn0
flabel comment s 4242 9043 4242 9043 0 FreeSans 800 0 0 0 dum
flabel comment s 5100 9043 5100 9043 0 FreeSans 800 0 0 0 Mn1
flabel comment s 5958 9043 5958 9043 0 FreeSans 800 0 0 0 Mn1
flabel comment s 6816 9043 6816 9043 0 FreeSans 800 0 0 0 dum
flabel metal2 9080 7636 9080 7636 0 FreeSans 1200 0 0 0 vbg_1v2
port 5 nsew
flabel metal1 8968 11290 8968 11290 0 FreeSans 800 0 0 0 vp
flabel metal3 9790 11203 9790 11203 0 FreeSans 1200 0 0 0 itest
port 2 nsew
flabel metal3 8074 11203 8074 11203 0 FreeSans 1200 0 0 0 ibias
port 3 nsew
flabel comment s 12820 10741 12820 10741 0 FreeSans 800 0 0 0 dum
flabel comment s 11962 10741 11962 10741 0 FreeSans 800 0 0 0 Mpp1
flabel comment s 11104 10741 11104 10741 0 FreeSans 800 0 0 0 Mpp1
flabel comment s 10246 10741 10246 10741 0 FreeSans 800 0 0 0 Mtst
flabel comment s 9388 10741 9388 10741 0 FreeSans 800 0 0 0 Mtst
flabel comment s 8530 10741 8530 10741 0 FreeSans 800 0 0 0 Mp
flabel comment s 7672 10741 7672 10741 0 FreeSans 800 0 0 0 Mp
flabel comment s 6814 10741 6814 10741 0 FreeSans 800 0 0 0 dum
flabel comment s 5956 10741 5956 10741 0 FreeSans 800 0 0 0 Mp1
flabel comment s 4240 10741 4240 10741 0 FreeSans 800 0 0 0 dum
flabel comment s 5098 10741 5098 10741 0 FreeSans 800 0 0 0 Mp1
flabel comment s 3382 10741 3382 10741 0 FreeSans 800 0 0 0 Mp0
flabel comment s 2524 10741 2524 10741 0 FreeSans 800 0 0 0 Mp0
flabel comment s 1666 10741 1666 10741 0 FreeSans 800 0 0 0 dum
flabel metal3 4674 10155 4674 10155 0 FreeSans 800 0 0 0 vp0
flabel space 10714 7425 10714 7425 0 FreeSans 480 0 0 0 M17
flabel space 10484 8834 10484 8834 0 FreeSans 480 0 0 0 Mt9
flabel space 11018 8834 11018 8834 0 FreeSans 480 0 0 0 Mt0
flabel space 11374 8834 11374 8834 0 FreeSans 480 0 0 0 Mt2
flabel metal3 10522 7346 10522 7346 0 FreeSans 800 0 0 0 vstart
flabel metal1 11197 8727 11197 8727 0 FreeSans 800 0 0 0 vp
flabel comment s 11737 8834 11737 8834 0 FreeSans 480 0 0 0 Mt7
flabel metal3 11626 8213 11626 8213 0 FreeSans 800 0 0 0 isrc_sel_b
flabel metal2 11723 7871 11723 7871 0 FreeSans 800 0 0 0 vn1
flabel metal3 11982 7648 11982 7648 0 FreeSans 1200 0 0 0 ena
port 7 nsew
flabel space 11148 636 11148 636 0 FreeSans 1600 0 0 0 Mnn1
flabel space 11148 1792 11148 1792 0 FreeSans 1600 0 0 0 Mnn1
flabel space 11148 4104 11148 4104 0 FreeSans 1600 0 0 0 Mnn1
flabel space 11148 5260 11148 5260 0 FreeSans 1600 0 0 0 Mnn1
flabel space 12806 5260 12806 5260 0 FreeSans 1600 0 0 0 Mnn1
flabel space 12806 4104 12806 4104 0 FreeSans 1600 0 0 0 Mnn1
flabel space 12806 2948 12806 2948 0 FreeSans 1600 0 0 0 Mnn0
flabel space 12806 1792 12806 1792 0 FreeSans 1600 0 0 0 Mnn1
flabel space 12806 636 12806 636 0 FreeSans 1600 0 0 0 Mnn1
flabel space 14464 636 14464 636 0 FreeSans 1600 0 0 0 dum
flabel space 14464 1792 14464 1792 0 FreeSans 1600 0 0 0 dum
flabel space 14464 2948 14464 2948 0 FreeSans 1600 0 0 0 dum
flabel space 14464 4104 14464 4104 0 FreeSans 1600 0 0 0 dum
flabel space 14464 5260 14464 5260 0 FreeSans 1600 0 0 0 dum
flabel space 9490 5260 9490 5260 0 FreeSans 1600 0 0 0 dum
flabel space 9490 4104 9490 4104 0 FreeSans 1600 0 0 0 dum
flabel space 9490 2948 9490 2948 0 FreeSans 1600 0 0 0 dum
flabel space 9490 1792 9490 1792 0 FreeSans 1600 0 0 0 dum
flabel space 9490 636 9490 636 0 FreeSans 1600 0 0 0 dum
flabel metal3 11786 7064 11786 7064 0 FreeSans 480 0 0 0 Mt6
flabel metal3 11964 7064 11964 7064 0 FreeSans 480 0 0 0 Mt4
flabel metal3 11602 7064 11602 7064 0 FreeSans 480 0 0 0 dum
flabel metal3 11424 7064 11424 7064 0 FreeSans 480 0 0 0 Mt3
flabel metal3 11246 7064 11246 7064 0 FreeSans 480 0 0 0 dum
flabel metal3 11068 7064 11068 7064 0 FreeSans 480 0 0 0 Mt1
flabel metal3 10890 7064 10890 7064 0 FreeSans 480 0 0 0 dum
flabel space 12720 7125 12720 7125 0 FreeSans 800 0 0 0 Ml9
flabel space 13178 7125 13178 7125 0 FreeSans 800 0 0 0 Ml10
flabel space 13636 7125 13636 7125 0 FreeSans 800 0 0 0 Ml1
flabel space 14094 7125 14094 7125 0 FreeSans 800 0 0 0 Ml0
flabel metal2 11517 7911 11517 7911 0 FreeSans 800 0 0 0 vp1
flabel metal3 1073 10722 1073 10722 0 FreeSans 1200 0 0 0 avdd
port 1 nsew
flabel comment s 10652 8834 10652 8834 0 FreeSans 480 0 0 0 Mt8
flabel comment s 10850 8836 10850 8836 0 FreeSans 480 0 0 0 dum
flabel comment s 11198 8834 11198 8836 0 FreeSans 480 0 0 0 dum
flabel comment s 11556 8834 11556 8834 0 FreeSans 480 0 0 0 dum
flabel comment s 11912 8836 11912 8836 0 FreeSans 480 0 0 0 Mt5
flabel space 12482 8848 12482 8848 0 FreeSans 800 0 0 0 Ml7
flabel space 12940 8848 12940 8848 0 FreeSans 800 0 0 0 Ml8
flabel space 13398 8848 13398 8848 0 FreeSans 800 0 0 0 Ml3
flabel space 13856 8848 13856 8848 0 FreeSans 800 0 0 0 Ml2
flabel space 14314 8848 14314 8848 0 FreeSans 800 0 0 0 Ml6
flabel metal2 s 13088 7824 13088 7824 0 FreeSans 800 0 0 0 ena_b
flabel comment s 14958 7108 14958 7108 0 FreeSans 800 0 0 0 Mn2
flabel comment s 15204 7104 15204 7104 0 FreeSans 800 0 0 0 dum
flabel comment s 15458 7083 15458 7083 0 FreeSans 800 0 0 0 Mn3
flabel comment s 14958 8813 14958 8813 0 FreeSans 800 0 0 0 Mp2
flabel comment s 15212 8809 15212 8809 0 FreeSans 800 0 0 0 dum
flabel comment s 15458 8809 15458 8809 0 FreeSans 800 0 0 0 Mp3
flabel metal3 10744 8129 10744 8129 0 FreeSans 1200 0 0 0 isrc_sel
port 6 nsew
flabel metal2 12034 8382 12034 8382 0 FreeSans 1200 0 0 0 ibg_200n
port 4 nsew
flabel metal3 s 3858 8771 3858 8771 0 FreeSans 1200 0 0 0 ve
port 9 nsew
<< end >>
