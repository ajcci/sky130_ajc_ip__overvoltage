magic
tech sky130A
magscale 1 2
timestamp 1711568248
<< nwell >>
rect -10177 -499 10177 499
<< mvpmos >>
rect -9919 118 -8319 202
rect -8261 118 -6661 202
rect -6603 118 -5003 202
rect -4945 118 -3345 202
rect -3287 118 -1687 202
rect -1629 118 -29 202
rect 29 118 1629 202
rect 1687 118 3287 202
rect 3345 118 4945 202
rect 5003 118 6603 202
rect 6661 118 8261 202
rect 8319 118 9919 202
rect -9919 -202 -8319 -118
rect -8261 -202 -6661 -118
rect -6603 -202 -5003 -118
rect -4945 -202 -3345 -118
rect -3287 -202 -1687 -118
rect -1629 -202 -29 -118
rect 29 -202 1629 -118
rect 1687 -202 3287 -118
rect 3345 -202 4945 -118
rect 5003 -202 6603 -118
rect 6661 -202 8261 -118
rect 8319 -202 9919 -118
<< mvpdiff >>
rect -9977 190 -9919 202
rect -9977 130 -9965 190
rect -9931 130 -9919 190
rect -9977 118 -9919 130
rect -8319 190 -8261 202
rect -8319 130 -8307 190
rect -8273 130 -8261 190
rect -8319 118 -8261 130
rect -6661 190 -6603 202
rect -6661 130 -6649 190
rect -6615 130 -6603 190
rect -6661 118 -6603 130
rect -5003 190 -4945 202
rect -5003 130 -4991 190
rect -4957 130 -4945 190
rect -5003 118 -4945 130
rect -3345 190 -3287 202
rect -3345 130 -3333 190
rect -3299 130 -3287 190
rect -3345 118 -3287 130
rect -1687 190 -1629 202
rect -1687 130 -1675 190
rect -1641 130 -1629 190
rect -1687 118 -1629 130
rect -29 190 29 202
rect -29 130 -17 190
rect 17 130 29 190
rect -29 118 29 130
rect 1629 190 1687 202
rect 1629 130 1641 190
rect 1675 130 1687 190
rect 1629 118 1687 130
rect 3287 190 3345 202
rect 3287 130 3299 190
rect 3333 130 3345 190
rect 3287 118 3345 130
rect 4945 190 5003 202
rect 4945 130 4957 190
rect 4991 130 5003 190
rect 4945 118 5003 130
rect 6603 190 6661 202
rect 6603 130 6615 190
rect 6649 130 6661 190
rect 6603 118 6661 130
rect 8261 190 8319 202
rect 8261 130 8273 190
rect 8307 130 8319 190
rect 8261 118 8319 130
rect 9919 190 9977 202
rect 9919 130 9931 190
rect 9965 130 9977 190
rect 9919 118 9977 130
rect -9977 -130 -9919 -118
rect -9977 -190 -9965 -130
rect -9931 -190 -9919 -130
rect -9977 -202 -9919 -190
rect -8319 -130 -8261 -118
rect -8319 -190 -8307 -130
rect -8273 -190 -8261 -130
rect -8319 -202 -8261 -190
rect -6661 -130 -6603 -118
rect -6661 -190 -6649 -130
rect -6615 -190 -6603 -130
rect -6661 -202 -6603 -190
rect -5003 -130 -4945 -118
rect -5003 -190 -4991 -130
rect -4957 -190 -4945 -130
rect -5003 -202 -4945 -190
rect -3345 -130 -3287 -118
rect -3345 -190 -3333 -130
rect -3299 -190 -3287 -130
rect -3345 -202 -3287 -190
rect -1687 -130 -1629 -118
rect -1687 -190 -1675 -130
rect -1641 -190 -1629 -130
rect -1687 -202 -1629 -190
rect -29 -130 29 -118
rect -29 -190 -17 -130
rect 17 -190 29 -130
rect -29 -202 29 -190
rect 1629 -130 1687 -118
rect 1629 -190 1641 -130
rect 1675 -190 1687 -130
rect 1629 -202 1687 -190
rect 3287 -130 3345 -118
rect 3287 -190 3299 -130
rect 3333 -190 3345 -130
rect 3287 -202 3345 -190
rect 4945 -130 5003 -118
rect 4945 -190 4957 -130
rect 4991 -190 5003 -130
rect 4945 -202 5003 -190
rect 6603 -130 6661 -118
rect 6603 -190 6615 -130
rect 6649 -190 6661 -130
rect 6603 -202 6661 -190
rect 8261 -130 8319 -118
rect 8261 -190 8273 -130
rect 8307 -190 8319 -130
rect 8261 -202 8319 -190
rect 9919 -130 9977 -118
rect 9919 -190 9931 -130
rect 9965 -190 9977 -130
rect 9919 -202 9977 -190
<< mvpdiffc >>
rect -9965 130 -9931 190
rect -8307 130 -8273 190
rect -6649 130 -6615 190
rect -4991 130 -4957 190
rect -3333 130 -3299 190
rect -1675 130 -1641 190
rect -17 130 17 190
rect 1641 130 1675 190
rect 3299 130 3333 190
rect 4957 130 4991 190
rect 6615 130 6649 190
rect 8273 130 8307 190
rect 9931 130 9965 190
rect -9965 -190 -9931 -130
rect -8307 -190 -8273 -130
rect -6649 -190 -6615 -130
rect -4991 -190 -4957 -130
rect -3333 -190 -3299 -130
rect -1675 -190 -1641 -130
rect -17 -190 17 -130
rect 1641 -190 1675 -130
rect 3299 -190 3333 -130
rect 4957 -190 4991 -130
rect 6615 -190 6649 -130
rect 8273 -190 8307 -130
rect 9931 -190 9965 -130
<< mvnsubdiff >>
rect -10111 421 10111 433
rect -10111 387 -10003 421
rect 10003 387 10111 421
rect -10111 375 10111 387
rect -10111 325 -10053 375
rect -10111 -325 -10099 325
rect -10065 -325 -10053 325
rect 10053 325 10111 375
rect -10111 -375 -10053 -325
rect 10053 -325 10065 325
rect 10099 -325 10111 325
rect 10053 -375 10111 -325
rect -10111 -387 10111 -375
rect -10111 -421 -10003 -387
rect 10003 -421 10111 -387
rect -10111 -433 10111 -421
<< mvnsubdiffcont >>
rect -10003 387 10003 421
rect -10099 -325 -10065 325
rect 10065 -325 10099 325
rect -10003 -421 10003 -387
<< poly >>
rect -9919 283 -8319 299
rect -9919 249 -9903 283
rect -8335 249 -8319 283
rect -9919 202 -8319 249
rect -8261 283 -6661 299
rect -8261 249 -8245 283
rect -6677 249 -6661 283
rect -8261 202 -6661 249
rect -6603 283 -5003 299
rect -6603 249 -6587 283
rect -5019 249 -5003 283
rect -6603 202 -5003 249
rect -4945 283 -3345 299
rect -4945 249 -4929 283
rect -3361 249 -3345 283
rect -4945 202 -3345 249
rect -3287 283 -1687 299
rect -3287 249 -3271 283
rect -1703 249 -1687 283
rect -3287 202 -1687 249
rect -1629 283 -29 299
rect -1629 249 -1613 283
rect -45 249 -29 283
rect -1629 202 -29 249
rect 29 283 1629 299
rect 29 249 45 283
rect 1613 249 1629 283
rect 29 202 1629 249
rect 1687 283 3287 299
rect 1687 249 1703 283
rect 3271 249 3287 283
rect 1687 202 3287 249
rect 3345 283 4945 299
rect 3345 249 3361 283
rect 4929 249 4945 283
rect 3345 202 4945 249
rect 5003 283 6603 299
rect 5003 249 5019 283
rect 6587 249 6603 283
rect 5003 202 6603 249
rect 6661 283 8261 299
rect 6661 249 6677 283
rect 8245 249 8261 283
rect 6661 202 8261 249
rect 8319 283 9919 299
rect 8319 249 8335 283
rect 9903 249 9919 283
rect 8319 202 9919 249
rect -9919 71 -8319 118
rect -9919 37 -9903 71
rect -8335 37 -8319 71
rect -9919 21 -8319 37
rect -8261 71 -6661 118
rect -8261 37 -8245 71
rect -6677 37 -6661 71
rect -8261 21 -6661 37
rect -6603 71 -5003 118
rect -6603 37 -6587 71
rect -5019 37 -5003 71
rect -6603 21 -5003 37
rect -4945 71 -3345 118
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -4945 21 -3345 37
rect -3287 71 -1687 118
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -3287 21 -1687 37
rect -1629 71 -29 118
rect -1629 37 -1613 71
rect -45 37 -29 71
rect -1629 21 -29 37
rect 29 71 1629 118
rect 29 37 45 71
rect 1613 37 1629 71
rect 29 21 1629 37
rect 1687 71 3287 118
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 1687 21 3287 37
rect 3345 71 4945 118
rect 3345 37 3361 71
rect 4929 37 4945 71
rect 3345 21 4945 37
rect 5003 71 6603 118
rect 5003 37 5019 71
rect 6587 37 6603 71
rect 5003 21 6603 37
rect 6661 71 8261 118
rect 6661 37 6677 71
rect 8245 37 8261 71
rect 6661 21 8261 37
rect 8319 71 9919 118
rect 8319 37 8335 71
rect 9903 37 9919 71
rect 8319 21 9919 37
rect -9919 -37 -8319 -21
rect -9919 -71 -9903 -37
rect -8335 -71 -8319 -37
rect -9919 -118 -8319 -71
rect -8261 -37 -6661 -21
rect -8261 -71 -8245 -37
rect -6677 -71 -6661 -37
rect -8261 -118 -6661 -71
rect -6603 -37 -5003 -21
rect -6603 -71 -6587 -37
rect -5019 -71 -5003 -37
rect -6603 -118 -5003 -71
rect -4945 -37 -3345 -21
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -4945 -118 -3345 -71
rect -3287 -37 -1687 -21
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -3287 -118 -1687 -71
rect -1629 -37 -29 -21
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect -1629 -118 -29 -71
rect 29 -37 1629 -21
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 29 -118 1629 -71
rect 1687 -37 3287 -21
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 1687 -118 3287 -71
rect 3345 -37 4945 -21
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect 3345 -118 4945 -71
rect 5003 -37 6603 -21
rect 5003 -71 5019 -37
rect 6587 -71 6603 -37
rect 5003 -118 6603 -71
rect 6661 -37 8261 -21
rect 6661 -71 6677 -37
rect 8245 -71 8261 -37
rect 6661 -118 8261 -71
rect 8319 -37 9919 -21
rect 8319 -71 8335 -37
rect 9903 -71 9919 -37
rect 8319 -118 9919 -71
rect -9919 -249 -8319 -202
rect -9919 -283 -9903 -249
rect -8335 -283 -8319 -249
rect -9919 -299 -8319 -283
rect -8261 -249 -6661 -202
rect -8261 -283 -8245 -249
rect -6677 -283 -6661 -249
rect -8261 -299 -6661 -283
rect -6603 -249 -5003 -202
rect -6603 -283 -6587 -249
rect -5019 -283 -5003 -249
rect -6603 -299 -5003 -283
rect -4945 -249 -3345 -202
rect -4945 -283 -4929 -249
rect -3361 -283 -3345 -249
rect -4945 -299 -3345 -283
rect -3287 -249 -1687 -202
rect -3287 -283 -3271 -249
rect -1703 -283 -1687 -249
rect -3287 -299 -1687 -283
rect -1629 -249 -29 -202
rect -1629 -283 -1613 -249
rect -45 -283 -29 -249
rect -1629 -299 -29 -283
rect 29 -249 1629 -202
rect 29 -283 45 -249
rect 1613 -283 1629 -249
rect 29 -299 1629 -283
rect 1687 -249 3287 -202
rect 1687 -283 1703 -249
rect 3271 -283 3287 -249
rect 1687 -299 3287 -283
rect 3345 -249 4945 -202
rect 3345 -283 3361 -249
rect 4929 -283 4945 -249
rect 3345 -299 4945 -283
rect 5003 -249 6603 -202
rect 5003 -283 5019 -249
rect 6587 -283 6603 -249
rect 5003 -299 6603 -283
rect 6661 -249 8261 -202
rect 6661 -283 6677 -249
rect 8245 -283 8261 -249
rect 6661 -299 8261 -283
rect 8319 -249 9919 -202
rect 8319 -283 8335 -249
rect 9903 -283 9919 -249
rect 8319 -299 9919 -283
<< polycont >>
rect -9903 249 -8335 283
rect -8245 249 -6677 283
rect -6587 249 -5019 283
rect -4929 249 -3361 283
rect -3271 249 -1703 283
rect -1613 249 -45 283
rect 45 249 1613 283
rect 1703 249 3271 283
rect 3361 249 4929 283
rect 5019 249 6587 283
rect 6677 249 8245 283
rect 8335 249 9903 283
rect -9903 37 -8335 71
rect -8245 37 -6677 71
rect -6587 37 -5019 71
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect 5019 37 6587 71
rect 6677 37 8245 71
rect 8335 37 9903 71
rect -9903 -71 -8335 -37
rect -8245 -71 -6677 -37
rect -6587 -71 -5019 -37
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
rect 5019 -71 6587 -37
rect 6677 -71 8245 -37
rect 8335 -71 9903 -37
rect -9903 -283 -8335 -249
rect -8245 -283 -6677 -249
rect -6587 -283 -5019 -249
rect -4929 -283 -3361 -249
rect -3271 -283 -1703 -249
rect -1613 -283 -45 -249
rect 45 -283 1613 -249
rect 1703 -283 3271 -249
rect 3361 -283 4929 -249
rect 5019 -283 6587 -249
rect 6677 -283 8245 -249
rect 8335 -283 9903 -249
<< locali >>
rect -10099 387 -10003 421
rect 10003 387 10099 421
rect -10099 325 -10065 387
rect 10065 325 10099 387
rect -9919 249 -9903 283
rect -8335 249 -8319 283
rect -8261 249 -8245 283
rect -6677 249 -6661 283
rect -6603 249 -6587 283
rect -5019 249 -5003 283
rect -4945 249 -4929 283
rect -3361 249 -3345 283
rect -3287 249 -3271 283
rect -1703 249 -1687 283
rect -1629 249 -1613 283
rect -45 249 -29 283
rect 29 249 45 283
rect 1613 249 1629 283
rect 1687 249 1703 283
rect 3271 249 3287 283
rect 3345 249 3361 283
rect 4929 249 4945 283
rect 5003 249 5019 283
rect 6587 249 6603 283
rect 6661 249 6677 283
rect 8245 249 8261 283
rect 8319 249 8335 283
rect 9903 249 9919 283
rect -9965 190 -9931 206
rect -9965 114 -9931 130
rect -8307 190 -8273 206
rect -8307 114 -8273 130
rect -6649 190 -6615 206
rect -6649 114 -6615 130
rect -4991 190 -4957 206
rect -4991 114 -4957 130
rect -3333 190 -3299 206
rect -3333 114 -3299 130
rect -1675 190 -1641 206
rect -1675 114 -1641 130
rect -17 190 17 206
rect -17 114 17 130
rect 1641 190 1675 206
rect 1641 114 1675 130
rect 3299 190 3333 206
rect 3299 114 3333 130
rect 4957 190 4991 206
rect 4957 114 4991 130
rect 6615 190 6649 206
rect 6615 114 6649 130
rect 8273 190 8307 206
rect 8273 114 8307 130
rect 9931 190 9965 206
rect 9931 114 9965 130
rect -9919 37 -9903 71
rect -8335 37 -8319 71
rect -8261 37 -8245 71
rect -6677 37 -6661 71
rect -6603 37 -6587 71
rect -5019 37 -5003 71
rect -4945 37 -4929 71
rect -3361 37 -3345 71
rect -3287 37 -3271 71
rect -1703 37 -1687 71
rect -1629 37 -1613 71
rect -45 37 -29 71
rect 29 37 45 71
rect 1613 37 1629 71
rect 1687 37 1703 71
rect 3271 37 3287 71
rect 3345 37 3361 71
rect 4929 37 4945 71
rect 5003 37 5019 71
rect 6587 37 6603 71
rect 6661 37 6677 71
rect 8245 37 8261 71
rect 8319 37 8335 71
rect 9903 37 9919 71
rect -9919 -71 -9903 -37
rect -8335 -71 -8319 -37
rect -8261 -71 -8245 -37
rect -6677 -71 -6661 -37
rect -6603 -71 -6587 -37
rect -5019 -71 -5003 -37
rect -4945 -71 -4929 -37
rect -3361 -71 -3345 -37
rect -3287 -71 -3271 -37
rect -1703 -71 -1687 -37
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 1687 -71 1703 -37
rect 3271 -71 3287 -37
rect 3345 -71 3361 -37
rect 4929 -71 4945 -37
rect 5003 -71 5019 -37
rect 6587 -71 6603 -37
rect 6661 -71 6677 -37
rect 8245 -71 8261 -37
rect 8319 -71 8335 -37
rect 9903 -71 9919 -37
rect -9965 -130 -9931 -114
rect -9965 -206 -9931 -190
rect -8307 -130 -8273 -114
rect -8307 -206 -8273 -190
rect -6649 -130 -6615 -114
rect -6649 -206 -6615 -190
rect -4991 -130 -4957 -114
rect -4991 -206 -4957 -190
rect -3333 -130 -3299 -114
rect -3333 -206 -3299 -190
rect -1675 -130 -1641 -114
rect -1675 -206 -1641 -190
rect -17 -130 17 -114
rect -17 -206 17 -190
rect 1641 -130 1675 -114
rect 1641 -206 1675 -190
rect 3299 -130 3333 -114
rect 3299 -206 3333 -190
rect 4957 -130 4991 -114
rect 4957 -206 4991 -190
rect 6615 -130 6649 -114
rect 6615 -206 6649 -190
rect 8273 -130 8307 -114
rect 8273 -206 8307 -190
rect 9931 -130 9965 -114
rect 9931 -206 9965 -190
rect -9919 -283 -9903 -249
rect -8335 -283 -8319 -249
rect -8261 -283 -8245 -249
rect -6677 -283 -6661 -249
rect -6603 -283 -6587 -249
rect -5019 -283 -5003 -249
rect -4945 -283 -4929 -249
rect -3361 -283 -3345 -249
rect -3287 -283 -3271 -249
rect -1703 -283 -1687 -249
rect -1629 -283 -1613 -249
rect -45 -283 -29 -249
rect 29 -283 45 -249
rect 1613 -283 1629 -249
rect 1687 -283 1703 -249
rect 3271 -283 3287 -249
rect 3345 -283 3361 -249
rect 4929 -283 4945 -249
rect 5003 -283 5019 -249
rect 6587 -283 6603 -249
rect 6661 -283 6677 -249
rect 8245 -283 8261 -249
rect 8319 -283 8335 -249
rect 9903 -283 9919 -249
rect -10099 -387 -10065 -325
rect 10065 -387 10099 -325
rect -10099 -421 -10003 -387
rect 10003 -421 10099 -387
<< viali >>
rect -9903 249 -8335 283
rect -8245 249 -6677 283
rect -6587 249 -5019 283
rect -4929 249 -3361 283
rect -3271 249 -1703 283
rect -1613 249 -45 283
rect 45 249 1613 283
rect 1703 249 3271 283
rect 3361 249 4929 283
rect 5019 249 6587 283
rect 6677 249 8245 283
rect 8335 249 9903 283
rect -9965 130 -9931 190
rect -8307 130 -8273 190
rect -6649 130 -6615 190
rect -4991 130 -4957 190
rect -3333 130 -3299 190
rect -1675 130 -1641 190
rect -17 130 17 190
rect 1641 130 1675 190
rect 3299 130 3333 190
rect 4957 130 4991 190
rect 6615 130 6649 190
rect 8273 130 8307 190
rect 9931 130 9965 190
rect -9903 37 -8335 71
rect -8245 37 -6677 71
rect -6587 37 -5019 71
rect -4929 37 -3361 71
rect -3271 37 -1703 71
rect -1613 37 -45 71
rect 45 37 1613 71
rect 1703 37 3271 71
rect 3361 37 4929 71
rect 5019 37 6587 71
rect 6677 37 8245 71
rect 8335 37 9903 71
rect -9903 -71 -8335 -37
rect -8245 -71 -6677 -37
rect -6587 -71 -5019 -37
rect -4929 -71 -3361 -37
rect -3271 -71 -1703 -37
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect 1703 -71 3271 -37
rect 3361 -71 4929 -37
rect 5019 -71 6587 -37
rect 6677 -71 8245 -37
rect 8335 -71 9903 -37
rect -9965 -190 -9931 -130
rect -8307 -190 -8273 -130
rect -6649 -190 -6615 -130
rect -4991 -190 -4957 -130
rect -3333 -190 -3299 -130
rect -1675 -190 -1641 -130
rect -17 -190 17 -130
rect 1641 -190 1675 -130
rect 3299 -190 3333 -130
rect 4957 -190 4991 -130
rect 6615 -190 6649 -130
rect 8273 -190 8307 -130
rect 9931 -190 9965 -130
rect -9903 -283 -8335 -249
rect -8245 -283 -6677 -249
rect -6587 -283 -5019 -249
rect -4929 -283 -3361 -249
rect -3271 -283 -1703 -249
rect -1613 -283 -45 -249
rect 45 -283 1613 -249
rect 1703 -283 3271 -249
rect 3361 -283 4929 -249
rect 5019 -283 6587 -249
rect 6677 -283 8245 -249
rect 8335 -283 9903 -249
<< metal1 >>
rect -9915 283 -8323 289
rect -9915 249 -9903 283
rect -8335 249 -8323 283
rect -9915 243 -8323 249
rect -8257 283 -6665 289
rect -8257 249 -8245 283
rect -6677 249 -6665 283
rect -8257 243 -6665 249
rect -6599 283 -5007 289
rect -6599 249 -6587 283
rect -5019 249 -5007 283
rect -6599 243 -5007 249
rect -4941 283 -3349 289
rect -4941 249 -4929 283
rect -3361 249 -3349 283
rect -4941 243 -3349 249
rect -3283 283 -1691 289
rect -3283 249 -3271 283
rect -1703 249 -1691 283
rect -3283 243 -1691 249
rect -1625 283 -33 289
rect -1625 249 -1613 283
rect -45 249 -33 283
rect -1625 243 -33 249
rect 33 283 1625 289
rect 33 249 45 283
rect 1613 249 1625 283
rect 33 243 1625 249
rect 1691 283 3283 289
rect 1691 249 1703 283
rect 3271 249 3283 283
rect 1691 243 3283 249
rect 3349 283 4941 289
rect 3349 249 3361 283
rect 4929 249 4941 283
rect 3349 243 4941 249
rect 5007 283 6599 289
rect 5007 249 5019 283
rect 6587 249 6599 283
rect 5007 243 6599 249
rect 6665 283 8257 289
rect 6665 249 6677 283
rect 8245 249 8257 283
rect 6665 243 8257 249
rect 8323 283 9915 289
rect 8323 249 8335 283
rect 9903 249 9915 283
rect 8323 243 9915 249
rect -9971 190 -9925 202
rect -9971 130 -9965 190
rect -9931 130 -9925 190
rect -9971 118 -9925 130
rect -8313 190 -8267 202
rect -8313 130 -8307 190
rect -8273 130 -8267 190
rect -8313 118 -8267 130
rect -6655 190 -6609 202
rect -6655 130 -6649 190
rect -6615 130 -6609 190
rect -6655 118 -6609 130
rect -4997 190 -4951 202
rect -4997 130 -4991 190
rect -4957 130 -4951 190
rect -4997 118 -4951 130
rect -3339 190 -3293 202
rect -3339 130 -3333 190
rect -3299 130 -3293 190
rect -3339 118 -3293 130
rect -1681 190 -1635 202
rect -1681 130 -1675 190
rect -1641 130 -1635 190
rect -1681 118 -1635 130
rect -23 190 23 202
rect -23 130 -17 190
rect 17 130 23 190
rect -23 118 23 130
rect 1635 190 1681 202
rect 1635 130 1641 190
rect 1675 130 1681 190
rect 1635 118 1681 130
rect 3293 190 3339 202
rect 3293 130 3299 190
rect 3333 130 3339 190
rect 3293 118 3339 130
rect 4951 190 4997 202
rect 4951 130 4957 190
rect 4991 130 4997 190
rect 4951 118 4997 130
rect 6609 190 6655 202
rect 6609 130 6615 190
rect 6649 130 6655 190
rect 6609 118 6655 130
rect 8267 190 8313 202
rect 8267 130 8273 190
rect 8307 130 8313 190
rect 8267 118 8313 130
rect 9925 190 9971 202
rect 9925 130 9931 190
rect 9965 130 9971 190
rect 9925 118 9971 130
rect -9915 71 -8323 77
rect -9915 37 -9903 71
rect -8335 37 -8323 71
rect -9915 31 -8323 37
rect -8257 71 -6665 77
rect -8257 37 -8245 71
rect -6677 37 -6665 71
rect -8257 31 -6665 37
rect -6599 71 -5007 77
rect -6599 37 -6587 71
rect -5019 37 -5007 71
rect -6599 31 -5007 37
rect -4941 71 -3349 77
rect -4941 37 -4929 71
rect -3361 37 -3349 71
rect -4941 31 -3349 37
rect -3283 71 -1691 77
rect -3283 37 -3271 71
rect -1703 37 -1691 71
rect -3283 31 -1691 37
rect -1625 71 -33 77
rect -1625 37 -1613 71
rect -45 37 -33 71
rect -1625 31 -33 37
rect 33 71 1625 77
rect 33 37 45 71
rect 1613 37 1625 71
rect 33 31 1625 37
rect 1691 71 3283 77
rect 1691 37 1703 71
rect 3271 37 3283 71
rect 1691 31 3283 37
rect 3349 71 4941 77
rect 3349 37 3361 71
rect 4929 37 4941 71
rect 3349 31 4941 37
rect 5007 71 6599 77
rect 5007 37 5019 71
rect 6587 37 6599 71
rect 5007 31 6599 37
rect 6665 71 8257 77
rect 6665 37 6677 71
rect 8245 37 8257 71
rect 6665 31 8257 37
rect 8323 71 9915 77
rect 8323 37 8335 71
rect 9903 37 9915 71
rect 8323 31 9915 37
rect -9915 -37 -8323 -31
rect -9915 -71 -9903 -37
rect -8335 -71 -8323 -37
rect -9915 -77 -8323 -71
rect -8257 -37 -6665 -31
rect -8257 -71 -8245 -37
rect -6677 -71 -6665 -37
rect -8257 -77 -6665 -71
rect -6599 -37 -5007 -31
rect -6599 -71 -6587 -37
rect -5019 -71 -5007 -37
rect -6599 -77 -5007 -71
rect -4941 -37 -3349 -31
rect -4941 -71 -4929 -37
rect -3361 -71 -3349 -37
rect -4941 -77 -3349 -71
rect -3283 -37 -1691 -31
rect -3283 -71 -3271 -37
rect -1703 -71 -1691 -37
rect -3283 -77 -1691 -71
rect -1625 -37 -33 -31
rect -1625 -71 -1613 -37
rect -45 -71 -33 -37
rect -1625 -77 -33 -71
rect 33 -37 1625 -31
rect 33 -71 45 -37
rect 1613 -71 1625 -37
rect 33 -77 1625 -71
rect 1691 -37 3283 -31
rect 1691 -71 1703 -37
rect 3271 -71 3283 -37
rect 1691 -77 3283 -71
rect 3349 -37 4941 -31
rect 3349 -71 3361 -37
rect 4929 -71 4941 -37
rect 3349 -77 4941 -71
rect 5007 -37 6599 -31
rect 5007 -71 5019 -37
rect 6587 -71 6599 -37
rect 5007 -77 6599 -71
rect 6665 -37 8257 -31
rect 6665 -71 6677 -37
rect 8245 -71 8257 -37
rect 6665 -77 8257 -71
rect 8323 -37 9915 -31
rect 8323 -71 8335 -37
rect 9903 -71 9915 -37
rect 8323 -77 9915 -71
rect -9971 -130 -9925 -118
rect -9971 -190 -9965 -130
rect -9931 -190 -9925 -130
rect -9971 -202 -9925 -190
rect -8313 -130 -8267 -118
rect -8313 -190 -8307 -130
rect -8273 -190 -8267 -130
rect -8313 -202 -8267 -190
rect -6655 -130 -6609 -118
rect -6655 -190 -6649 -130
rect -6615 -190 -6609 -130
rect -6655 -202 -6609 -190
rect -4997 -130 -4951 -118
rect -4997 -190 -4991 -130
rect -4957 -190 -4951 -130
rect -4997 -202 -4951 -190
rect -3339 -130 -3293 -118
rect -3339 -190 -3333 -130
rect -3299 -190 -3293 -130
rect -3339 -202 -3293 -190
rect -1681 -130 -1635 -118
rect -1681 -190 -1675 -130
rect -1641 -190 -1635 -130
rect -1681 -202 -1635 -190
rect -23 -130 23 -118
rect -23 -190 -17 -130
rect 17 -190 23 -130
rect -23 -202 23 -190
rect 1635 -130 1681 -118
rect 1635 -190 1641 -130
rect 1675 -190 1681 -130
rect 1635 -202 1681 -190
rect 3293 -130 3339 -118
rect 3293 -190 3299 -130
rect 3333 -190 3339 -130
rect 3293 -202 3339 -190
rect 4951 -130 4997 -118
rect 4951 -190 4957 -130
rect 4991 -190 4997 -130
rect 4951 -202 4997 -190
rect 6609 -130 6655 -118
rect 6609 -190 6615 -130
rect 6649 -190 6655 -130
rect 6609 -202 6655 -190
rect 8267 -130 8313 -118
rect 8267 -190 8273 -130
rect 8307 -190 8313 -130
rect 8267 -202 8313 -190
rect 9925 -130 9971 -118
rect 9925 -190 9931 -130
rect 9965 -190 9971 -130
rect 9925 -202 9971 -190
rect -9915 -249 -8323 -243
rect -9915 -283 -9903 -249
rect -8335 -283 -8323 -249
rect -9915 -289 -8323 -283
rect -8257 -249 -6665 -243
rect -8257 -283 -8245 -249
rect -6677 -283 -6665 -249
rect -8257 -289 -6665 -283
rect -6599 -249 -5007 -243
rect -6599 -283 -6587 -249
rect -5019 -283 -5007 -249
rect -6599 -289 -5007 -283
rect -4941 -249 -3349 -243
rect -4941 -283 -4929 -249
rect -3361 -283 -3349 -249
rect -4941 -289 -3349 -283
rect -3283 -249 -1691 -243
rect -3283 -283 -3271 -249
rect -1703 -283 -1691 -249
rect -3283 -289 -1691 -283
rect -1625 -249 -33 -243
rect -1625 -283 -1613 -249
rect -45 -283 -33 -249
rect -1625 -289 -33 -283
rect 33 -249 1625 -243
rect 33 -283 45 -249
rect 1613 -283 1625 -249
rect 33 -289 1625 -283
rect 1691 -249 3283 -243
rect 1691 -283 1703 -249
rect 3271 -283 3283 -249
rect 1691 -289 3283 -283
rect 3349 -249 4941 -243
rect 3349 -283 3361 -249
rect 4929 -283 4941 -249
rect 3349 -289 4941 -283
rect 5007 -249 6599 -243
rect 5007 -283 5019 -249
rect 6587 -283 6599 -249
rect 5007 -289 6599 -283
rect 6665 -249 8257 -243
rect 6665 -283 6677 -249
rect 8245 -283 8257 -249
rect 6665 -289 8257 -283
rect 8323 -249 9915 -243
rect 8323 -283 8335 -249
rect 9903 -283 9915 -249
rect 8323 -289 9915 -283
<< properties >>
string FIXED_BBOX -10082 -404 10082 404
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 8.0 m 2 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
