magic
tech sky130A
magscale 1 2
timestamp 1711636687
<< nwell >>
rect -407 -347 407 347
<< mvpmos >>
rect -149 -50 -29 50
rect 29 -50 149 50
<< mvpdiff >>
rect -207 38 -149 50
rect -207 -38 -195 38
rect -161 -38 -149 38
rect -207 -50 -149 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 149 38 207 50
rect 149 -38 161 38
rect 195 -38 207 38
rect 149 -50 207 -38
<< mvpdiffc >>
rect -195 -38 -161 38
rect -17 -38 17 38
rect 161 -38 195 38
<< mvnsubdiff >>
rect -341 269 341 281
rect -341 235 -233 269
rect 233 235 341 269
rect -341 223 341 235
rect -341 173 -283 223
rect -341 -173 -329 173
rect -295 -173 -283 173
rect 283 173 341 223
rect -341 -223 -283 -173
rect 283 -173 295 173
rect 329 -173 341 173
rect 283 -223 341 -173
rect -341 -235 341 -223
rect -341 -269 -233 -235
rect 233 -269 341 -235
rect -341 -281 341 -269
<< mvnsubdiffcont >>
rect -233 235 233 269
rect -329 -173 -295 173
rect 295 -173 329 173
rect -233 -269 233 -235
<< poly >>
rect -149 131 -29 147
rect -149 97 -133 131
rect -45 97 -29 131
rect -149 50 -29 97
rect 29 131 149 147
rect 29 97 45 131
rect 133 97 149 131
rect 29 50 149 97
rect -149 -97 -29 -50
rect -149 -131 -133 -97
rect -45 -131 -29 -97
rect -149 -147 -29 -131
rect 29 -97 149 -50
rect 29 -131 45 -97
rect 133 -131 149 -97
rect 29 -147 149 -131
<< polycont >>
rect -133 97 -45 131
rect 45 97 133 131
rect -133 -131 -45 -97
rect 45 -131 133 -97
<< locali >>
rect -329 235 -233 269
rect 233 235 329 269
rect -329 173 -295 235
rect 295 173 329 235
rect -149 97 -133 131
rect -45 97 -29 131
rect 29 97 45 131
rect 133 97 149 131
rect -195 38 -161 54
rect -195 -54 -161 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 161 38 195 54
rect 161 -54 195 -38
rect -149 -131 -133 -97
rect -45 -131 -29 -97
rect 29 -131 45 -97
rect 133 -131 149 -97
rect -329 -235 -295 -173
rect 295 -235 329 -173
rect -329 -269 -233 -235
rect 233 -269 329 -235
<< viali >>
rect -133 97 -45 131
rect 45 97 133 131
rect -195 -38 -161 38
rect -17 -38 17 38
rect 161 -38 195 38
rect -133 -131 -45 -97
rect 45 -131 133 -97
<< metal1 >>
rect -145 131 -33 137
rect -145 97 -133 131
rect -45 97 -33 131
rect -145 91 -33 97
rect 33 131 145 137
rect 33 97 45 131
rect 133 97 145 131
rect 33 91 145 97
rect -201 38 -155 50
rect -201 -38 -195 38
rect -161 -38 -155 38
rect -201 -50 -155 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 155 38 201 50
rect 155 -38 161 38
rect 195 -38 201 38
rect 155 -50 201 -38
rect -145 -97 -33 -91
rect -145 -131 -133 -97
rect -45 -131 -33 -97
rect -145 -137 -33 -131
rect 33 -97 145 -91
rect 33 -131 45 -97
rect 133 -131 145 -97
rect 33 -137 145 -131
<< properties >>
string FIXED_BBOX -312 -252 312 252
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 0.6 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
