* NGSPICE file created from overvoltage_dig.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
X0 Y a_91_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_91_199# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_341_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X6 a_245_297# C a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7 a_341_297# B a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X8 a_91_199# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X9 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.52 ps=3.04 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt overvoltage_dig VPWR otrip_decoded[15] otrip_decoded[14] otrip_decoded[13]
+ otrip_decoded[12] otrip_decoded[11] otrip_decoded[10] otrip_decoded[9] otrip_decoded[8]
+ otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[4] otrip_decoded[3]
+ otrip_decoded[2] otrip_decoded[1] otrip_decoded[0] VGND otrip[3] otrip[2] otrip[1]
+ otrip[0]
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput20 net20 VGND VGND VPWR VPWR otrip_decoded[9] sky130_fd_sc_hd__buf_2
Xoutput7 net7 VGND VGND VPWR VPWR otrip_decoded[11] sky130_fd_sc_hd__buf_2
XFILLER_0_13_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput10 net10 VGND VGND VPWR VPWR otrip_decoded[14] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput8 net8 VGND VGND VPWR VPWR otrip_decoded[12] sky130_fd_sc_hd__buf_2
XFILLER_0_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR otrip_decoded[13] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR otrip_decoded[15] sky130_fd_sc_hd__buf_2
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__buf_2
XFILLER_0_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput13 net13 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_4_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__buf_2
X_09_ net25 net23 net22 net28 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08_ net28 net26 net24 net22 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__nor4b_1
XFILLER_0_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__buf_2
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07_ net21 net27 net26 net24 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__and4b_1
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__buf_2
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__buf_2
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06_ net21 net27 net25 net23 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__and4bb_1
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput19 net19 VGND VGND VPWR VPWR otrip_decoded[8] sky130_fd_sc_hd__buf_2
X_05_ net21 net25 net23 net27 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__and4bb_1
XFILLER_0_13_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout21 net4 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04_ net21 net27 net25 net23 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__nor4b_1
XFILLER_0_2_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout22 net4 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput1 otrip[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_03_ net21 net23 net25 net27 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout23 net3 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 otrip[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_3_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_02_ net21 net27 net23 net25 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor4b_1
XFILLER_0_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout24 net3 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
X_01_ net21 net25 net23 net27 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__nor4b_1
Xinput3 otrip[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout25 net2 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 otrip[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_00_ net21 net27 net25 net23 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__nor4_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout26 net2 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout27 net1 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout28 net1 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_11 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15_ net22 net28 net26 net24 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__and4_1
XFILLER_0_0_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14_ net28 net26 net24 net22 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__and4b_1
XFILLER_0_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13_ net26 net24 net22 net28 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12_ net27 net25 net23 net21 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11_ net24 net26 net28 net22 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__and4b_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10_ net27 net23 net25 net21 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput5 net5 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__buf_2
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput6 net6 VGND VGND VPWR VPWR otrip_decoded[10] sky130_fd_sc_hd__buf_2
.ends

