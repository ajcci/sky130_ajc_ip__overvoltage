magic
tech sky130A
magscale 1 2
timestamp 1711690227
<< pwell >>
rect 19634 -5518 20560 -4674
<< mvnmos >>
rect 19985 -5183 20085 -5099
<< mvndiff >>
rect 19927 -5111 19985 -5099
rect 19927 -5171 19939 -5111
rect 19973 -5171 19985 -5111
rect 19927 -5183 19985 -5171
rect 20085 -5111 20143 -5099
rect 20085 -5171 20097 -5111
rect 20131 -5171 20143 -5111
rect 20085 -5183 20143 -5171
<< mvndiffc >>
rect 19939 -5171 19973 -5111
rect 20097 -5171 20131 -5111
<< mvpsubdiff >>
rect 20278 -4904 20384 -4802
rect 20278 -4924 20344 -4904
rect 20362 -4924 20384 -4904
rect 20278 -4998 20384 -4924
<< mvpsubdiffcont >>
rect 20344 -4924 20362 -4904
<< poly >>
rect 19985 -5027 20085 -5011
rect 19985 -5061 20001 -5027
rect 20069 -5061 20085 -5027
rect 19985 -5099 20085 -5061
rect 19985 -5221 20085 -5183
rect 19985 -5255 20001 -5221
rect 20069 -5255 20085 -5221
rect 19985 -5271 20085 -5255
<< polycont >>
rect 20001 -5061 20069 -5027
rect 20001 -5255 20069 -5221
<< locali >>
rect 20248 -4904 20403 -4889
rect 20248 -4924 20344 -4904
rect 20362 -4924 20403 -4904
rect 20248 -4936 20403 -4924
rect 19985 -5061 20001 -5027
rect 20069 -5061 20085 -5027
rect 19939 -5111 19973 -5095
rect 19939 -5187 19973 -5171
rect 20097 -5111 20131 -5095
rect 20097 -5187 20131 -5171
rect 19985 -5255 20001 -5221
rect 20069 -5255 20085 -5221
<< viali >>
rect 20001 -5061 20069 -5027
rect 19939 -5171 19973 -5111
rect 20097 -5171 20131 -5111
rect 20001 -5255 20069 -5221
<< metal1 >>
rect 19985 -5027 20081 -5021
rect 19985 -5061 20001 -5027
rect 20069 -5061 20081 -5027
rect 19985 -5067 20081 -5061
rect 19933 -5111 19979 -5095
rect 19933 -5171 19939 -5111
rect 19973 -5171 19979 -5111
rect 19933 -5183 19979 -5171
rect 20091 -5111 20137 -5095
rect 20091 -5171 20097 -5111
rect 20131 -5171 20137 -5111
rect 20091 -5183 20137 -5171
rect 19989 -5221 20081 -5215
rect 19989 -5255 20001 -5221
rect 20069 -5255 20081 -5221
rect 19989 -5261 20081 -5255
<< end >>
