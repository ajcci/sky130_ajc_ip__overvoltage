magic
tech sky130A
magscale 1 2
timestamp 1712109191
<< pwell >>
rect -3515 -3039 3515 3039
<< mvnmos >>
rect -3287 1781 -1687 2781
rect -1629 1781 -29 2781
rect 29 1781 1629 2781
rect 1687 1781 3287 2781
rect -3287 625 -1687 1625
rect -1629 625 -29 1625
rect 29 625 1629 1625
rect 1687 625 3287 1625
rect -3287 -531 -1687 469
rect -1629 -531 -29 469
rect 29 -531 1629 469
rect 1687 -531 3287 469
rect -3287 -1687 -1687 -687
rect -1629 -1687 -29 -687
rect 29 -1687 1629 -687
rect 1687 -1687 3287 -687
rect -3287 -2843 -1687 -1843
rect -1629 -2843 -29 -1843
rect 29 -2843 1629 -1843
rect 1687 -2843 3287 -1843
<< mvndiff >>
rect -3345 2769 -3287 2781
rect -3345 1793 -3333 2769
rect -3299 1793 -3287 2769
rect -3345 1781 -3287 1793
rect -1687 2769 -1629 2781
rect -1687 1793 -1675 2769
rect -1641 1793 -1629 2769
rect -1687 1781 -1629 1793
rect -29 2769 29 2781
rect -29 1793 -17 2769
rect 17 1793 29 2769
rect -29 1781 29 1793
rect 1629 2769 1687 2781
rect 1629 1793 1641 2769
rect 1675 1793 1687 2769
rect 1629 1781 1687 1793
rect 3287 2769 3345 2781
rect 3287 1793 3299 2769
rect 3333 1793 3345 2769
rect 3287 1781 3345 1793
rect -3345 1613 -3287 1625
rect -3345 637 -3333 1613
rect -3299 637 -3287 1613
rect -3345 625 -3287 637
rect -1687 1613 -1629 1625
rect -1687 637 -1675 1613
rect -1641 637 -1629 1613
rect -1687 625 -1629 637
rect -29 1613 29 1625
rect -29 637 -17 1613
rect 17 637 29 1613
rect -29 625 29 637
rect 1629 1613 1687 1625
rect 1629 637 1641 1613
rect 1675 637 1687 1613
rect 1629 625 1687 637
rect 3287 1613 3345 1625
rect 3287 637 3299 1613
rect 3333 637 3345 1613
rect 3287 625 3345 637
rect -3345 457 -3287 469
rect -3345 -519 -3333 457
rect -3299 -519 -3287 457
rect -3345 -531 -3287 -519
rect -1687 457 -1629 469
rect -1687 -519 -1675 457
rect -1641 -519 -1629 457
rect -1687 -531 -1629 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 1629 457 1687 469
rect 1629 -519 1641 457
rect 1675 -519 1687 457
rect 1629 -531 1687 -519
rect 3287 457 3345 469
rect 3287 -519 3299 457
rect 3333 -519 3345 457
rect 3287 -531 3345 -519
rect -3345 -699 -3287 -687
rect -3345 -1675 -3333 -699
rect -3299 -1675 -3287 -699
rect -3345 -1687 -3287 -1675
rect -1687 -699 -1629 -687
rect -1687 -1675 -1675 -699
rect -1641 -1675 -1629 -699
rect -1687 -1687 -1629 -1675
rect -29 -699 29 -687
rect -29 -1675 -17 -699
rect 17 -1675 29 -699
rect -29 -1687 29 -1675
rect 1629 -699 1687 -687
rect 1629 -1675 1641 -699
rect 1675 -1675 1687 -699
rect 1629 -1687 1687 -1675
rect 3287 -699 3345 -687
rect 3287 -1675 3299 -699
rect 3333 -1675 3345 -699
rect 3287 -1687 3345 -1675
rect -3345 -1855 -3287 -1843
rect -3345 -2831 -3333 -1855
rect -3299 -2831 -3287 -1855
rect -3345 -2843 -3287 -2831
rect -1687 -1855 -1629 -1843
rect -1687 -2831 -1675 -1855
rect -1641 -2831 -1629 -1855
rect -1687 -2843 -1629 -2831
rect -29 -1855 29 -1843
rect -29 -2831 -17 -1855
rect 17 -2831 29 -1855
rect -29 -2843 29 -2831
rect 1629 -1855 1687 -1843
rect 1629 -2831 1641 -1855
rect 1675 -2831 1687 -1855
rect 1629 -2843 1687 -2831
rect 3287 -1855 3345 -1843
rect 3287 -2831 3299 -1855
rect 3333 -2831 3345 -1855
rect 3287 -2843 3345 -2831
<< mvndiffc >>
rect -3333 1793 -3299 2769
rect -1675 1793 -1641 2769
rect -17 1793 17 2769
rect 1641 1793 1675 2769
rect 3299 1793 3333 2769
rect -3333 637 -3299 1613
rect -1675 637 -1641 1613
rect -17 637 17 1613
rect 1641 637 1675 1613
rect 3299 637 3333 1613
rect -3333 -519 -3299 457
rect -1675 -519 -1641 457
rect -17 -519 17 457
rect 1641 -519 1675 457
rect 3299 -519 3333 457
rect -3333 -1675 -3299 -699
rect -1675 -1675 -1641 -699
rect -17 -1675 17 -699
rect 1641 -1675 1675 -699
rect 3299 -1675 3333 -699
rect -3333 -2831 -3299 -1855
rect -1675 -2831 -1641 -1855
rect -17 -2831 17 -1855
rect 1641 -2831 1675 -1855
rect 3299 -2831 3333 -1855
<< mvpsubdiff >>
rect -3479 2991 3479 3003
rect -3479 2957 -3371 2991
rect 3371 2957 3479 2991
rect -3479 2945 3479 2957
rect -3479 2895 -3421 2945
rect -3479 -2895 -3467 2895
rect -3433 -2895 -3421 2895
rect 3421 2895 3479 2945
rect -3479 -2945 -3421 -2895
rect 3421 -2895 3433 2895
rect 3467 -2895 3479 2895
rect 3421 -2945 3479 -2895
rect -3479 -2957 3479 -2945
rect -3479 -2991 -3371 -2957
rect 3371 -2991 3479 -2957
rect -3479 -3003 3479 -2991
<< mvpsubdiffcont >>
rect -3371 2957 3371 2991
rect -3467 -2895 -3433 2895
rect 3433 -2895 3467 2895
rect -3371 -2991 3371 -2957
<< poly >>
rect -3287 2853 -1687 2869
rect -3287 2819 -3271 2853
rect -1703 2819 -1687 2853
rect -3287 2781 -1687 2819
rect -1629 2853 -29 2869
rect -1629 2819 -1613 2853
rect -45 2819 -29 2853
rect -1629 2781 -29 2819
rect 29 2853 1629 2869
rect 29 2819 45 2853
rect 1613 2819 1629 2853
rect 29 2781 1629 2819
rect 1687 2853 3287 2869
rect 1687 2819 1703 2853
rect 3271 2819 3287 2853
rect 1687 2781 3287 2819
rect -3287 1755 -1687 1781
rect -1629 1755 -29 1781
rect 29 1755 1629 1781
rect 1687 1755 3287 1781
rect -3287 1697 -1687 1713
rect -3287 1663 -3271 1697
rect -1703 1663 -1687 1697
rect -3287 1625 -1687 1663
rect -1629 1697 -29 1713
rect -1629 1663 -1613 1697
rect -45 1663 -29 1697
rect -1629 1625 -29 1663
rect 29 1697 1629 1713
rect 29 1663 45 1697
rect 1613 1663 1629 1697
rect 29 1625 1629 1663
rect 1687 1697 3287 1713
rect 1687 1663 1703 1697
rect 3271 1663 3287 1697
rect 1687 1625 3287 1663
rect -3287 599 -1687 625
rect -1629 599 -29 625
rect 29 599 1629 625
rect 1687 599 3287 625
rect -3287 541 -1687 557
rect -3287 507 -3271 541
rect -1703 507 -1687 541
rect -3287 469 -1687 507
rect -1629 541 -29 557
rect -1629 507 -1613 541
rect -45 507 -29 541
rect -1629 469 -29 507
rect 29 541 1629 557
rect 29 507 45 541
rect 1613 507 1629 541
rect 29 469 1629 507
rect 1687 541 3287 557
rect 1687 507 1703 541
rect 3271 507 3287 541
rect 1687 469 3287 507
rect -3287 -557 -1687 -531
rect -1629 -557 -29 -531
rect 29 -557 1629 -531
rect 1687 -557 3287 -531
rect -3287 -615 -1687 -599
rect -3287 -649 -3271 -615
rect -1703 -649 -1687 -615
rect -3287 -687 -1687 -649
rect -1629 -615 -29 -599
rect -1629 -649 -1613 -615
rect -45 -649 -29 -615
rect -1629 -687 -29 -649
rect 29 -615 1629 -599
rect 29 -649 45 -615
rect 1613 -649 1629 -615
rect 29 -687 1629 -649
rect 1687 -615 3287 -599
rect 1687 -649 1703 -615
rect 3271 -649 3287 -615
rect 1687 -687 3287 -649
rect -3287 -1713 -1687 -1687
rect -1629 -1713 -29 -1687
rect 29 -1713 1629 -1687
rect 1687 -1713 3287 -1687
rect -3287 -1771 -1687 -1755
rect -3287 -1805 -3271 -1771
rect -1703 -1805 -1687 -1771
rect -3287 -1843 -1687 -1805
rect -1629 -1771 -29 -1755
rect -1629 -1805 -1613 -1771
rect -45 -1805 -29 -1771
rect -1629 -1843 -29 -1805
rect 29 -1771 1629 -1755
rect 29 -1805 45 -1771
rect 1613 -1805 1629 -1771
rect 29 -1843 1629 -1805
rect 1687 -1771 3287 -1755
rect 1687 -1805 1703 -1771
rect 3271 -1805 3287 -1771
rect 1687 -1843 3287 -1805
rect -3287 -2869 -1687 -2843
rect -1629 -2869 -29 -2843
rect 29 -2869 1629 -2843
rect 1687 -2869 3287 -2843
<< polycont >>
rect -3271 2819 -1703 2853
rect -1613 2819 -45 2853
rect 45 2819 1613 2853
rect 1703 2819 3271 2853
rect -3271 1663 -1703 1697
rect -1613 1663 -45 1697
rect 45 1663 1613 1697
rect 1703 1663 3271 1697
rect -3271 507 -1703 541
rect -1613 507 -45 541
rect 45 507 1613 541
rect 1703 507 3271 541
rect -3271 -649 -1703 -615
rect -1613 -649 -45 -615
rect 45 -649 1613 -615
rect 1703 -649 3271 -615
rect -3271 -1805 -1703 -1771
rect -1613 -1805 -45 -1771
rect 45 -1805 1613 -1771
rect 1703 -1805 3271 -1771
<< locali >>
rect -3467 2957 -3371 2991
rect 3371 2957 3467 2991
rect -3467 2895 -3433 2957
rect 3433 2895 3467 2957
rect -3287 2819 -3271 2853
rect -1703 2819 -1687 2853
rect -1629 2819 -1613 2853
rect -45 2819 -29 2853
rect 29 2819 45 2853
rect 1613 2819 1629 2853
rect 1687 2819 1703 2853
rect 3271 2819 3287 2853
rect -3333 2769 -3299 2785
rect -3333 1777 -3299 1793
rect -1675 2769 -1641 2785
rect -1675 1777 -1641 1793
rect -17 2769 17 2785
rect -17 1777 17 1793
rect 1641 2769 1675 2785
rect 1641 1777 1675 1793
rect 3299 2769 3333 2785
rect 3299 1777 3333 1793
rect -3287 1663 -3271 1697
rect -1703 1663 -1687 1697
rect -1629 1663 -1613 1697
rect -45 1663 -29 1697
rect 29 1663 45 1697
rect 1613 1663 1629 1697
rect 1687 1663 1703 1697
rect 3271 1663 3287 1697
rect -3333 1613 -3299 1629
rect -3333 621 -3299 637
rect -1675 1613 -1641 1629
rect -1675 621 -1641 637
rect -17 1613 17 1629
rect -17 621 17 637
rect 1641 1613 1675 1629
rect 1641 621 1675 637
rect 3299 1613 3333 1629
rect 3299 621 3333 637
rect -3287 507 -3271 541
rect -1703 507 -1687 541
rect -1629 507 -1613 541
rect -45 507 -29 541
rect 29 507 45 541
rect 1613 507 1629 541
rect 1687 507 1703 541
rect 3271 507 3287 541
rect -3333 457 -3299 473
rect -3333 -535 -3299 -519
rect -1675 457 -1641 473
rect -1675 -535 -1641 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 1641 457 1675 473
rect 1641 -535 1675 -519
rect 3299 457 3333 473
rect 3299 -535 3333 -519
rect -3287 -649 -3271 -615
rect -1703 -649 -1687 -615
rect -1629 -649 -1613 -615
rect -45 -649 -29 -615
rect 29 -649 45 -615
rect 1613 -649 1629 -615
rect 1687 -649 1703 -615
rect 3271 -649 3287 -615
rect -3333 -699 -3299 -683
rect -3333 -1691 -3299 -1675
rect -1675 -699 -1641 -683
rect -1675 -1691 -1641 -1675
rect -17 -699 17 -683
rect -17 -1691 17 -1675
rect 1641 -699 1675 -683
rect 1641 -1691 1675 -1675
rect 3299 -699 3333 -683
rect 3299 -1691 3333 -1675
rect -3287 -1805 -3271 -1771
rect -1703 -1805 -1687 -1771
rect -1629 -1805 -1613 -1771
rect -45 -1805 -29 -1771
rect 29 -1805 45 -1771
rect 1613 -1805 1629 -1771
rect 1687 -1805 1703 -1771
rect 3271 -1805 3287 -1771
rect -3333 -1855 -3299 -1839
rect -3333 -2847 -3299 -2831
rect -1675 -1855 -1641 -1839
rect -1675 -2847 -1641 -2831
rect -17 -1855 17 -1839
rect -17 -2847 17 -2831
rect 1641 -1855 1675 -1839
rect 1641 -2847 1675 -2831
rect 3299 -1855 3333 -1839
rect 3299 -2847 3333 -2831
rect -3467 -2957 -3433 -2895
rect 3433 -2957 3467 -2895
rect -3467 -2991 -3371 -2957
rect 3371 -2991 3467 -2957
<< viali >>
rect -3271 2819 -1703 2853
rect -1613 2819 -45 2853
rect 45 2819 1613 2853
rect 1703 2819 3271 2853
rect -3333 1793 -3299 2769
rect -1675 1793 -1641 2769
rect -17 1793 17 2769
rect 1641 1793 1675 2769
rect 3299 1793 3333 2769
rect -3271 1663 -1703 1697
rect -1613 1663 -45 1697
rect 45 1663 1613 1697
rect 1703 1663 3271 1697
rect -3333 637 -3299 1613
rect -1675 637 -1641 1613
rect -17 637 17 1613
rect 1641 637 1675 1613
rect 3299 637 3333 1613
rect -3271 507 -1703 541
rect -1613 507 -45 541
rect 45 507 1613 541
rect 1703 507 3271 541
rect -3333 -519 -3299 457
rect -1675 -519 -1641 457
rect -17 -519 17 457
rect 1641 -519 1675 457
rect 3299 -519 3333 457
rect -3271 -649 -1703 -615
rect -1613 -649 -45 -615
rect 45 -649 1613 -615
rect 1703 -649 3271 -615
rect -3333 -1675 -3299 -699
rect -1675 -1675 -1641 -699
rect -17 -1675 17 -699
rect 1641 -1675 1675 -699
rect 3299 -1675 3333 -699
rect -3271 -1805 -1703 -1771
rect -1613 -1805 -45 -1771
rect 45 -1805 1613 -1771
rect 1703 -1805 3271 -1771
rect -3333 -2831 -3299 -1855
rect -1675 -2831 -1641 -1855
rect -17 -2831 17 -1855
rect 1641 -2831 1675 -1855
rect 3299 -2831 3333 -1855
<< metal1 >>
rect -3283 2853 -1691 2859
rect -3283 2819 -3271 2853
rect -1703 2819 -1691 2853
rect -3283 2813 -1691 2819
rect -1625 2853 -33 2859
rect -1625 2819 -1613 2853
rect -45 2819 -33 2853
rect -1625 2813 -33 2819
rect 33 2853 1625 2859
rect 33 2819 45 2853
rect 1613 2819 1625 2853
rect 33 2813 1625 2819
rect 1691 2853 3283 2859
rect 1691 2819 1703 2853
rect 3271 2819 3283 2853
rect 1691 2813 3283 2819
rect -3339 2769 -3293 2781
rect -3339 1793 -3333 2769
rect -3299 1793 -3293 2769
rect -3339 1781 -3293 1793
rect -1681 2769 -1635 2781
rect -1681 1793 -1675 2769
rect -1641 1793 -1635 2769
rect -1681 1781 -1635 1793
rect -23 2769 23 2781
rect -23 1793 -17 2769
rect 17 1793 23 2769
rect -23 1781 23 1793
rect 1635 2769 1681 2781
rect 1635 1793 1641 2769
rect 1675 1793 1681 2769
rect 1635 1781 1681 1793
rect 3293 2769 3339 2781
rect 3293 1793 3299 2769
rect 3333 1793 3339 2769
rect 3293 1781 3339 1793
rect -3283 1697 -1691 1703
rect -3283 1663 -3271 1697
rect -1703 1663 -1691 1697
rect -3283 1657 -1691 1663
rect -1625 1697 -33 1703
rect -1625 1663 -1613 1697
rect -45 1663 -33 1697
rect -1625 1657 -33 1663
rect 33 1697 1625 1703
rect 33 1663 45 1697
rect 1613 1663 1625 1697
rect 33 1657 1625 1663
rect 1691 1697 3283 1703
rect 1691 1663 1703 1697
rect 3271 1663 3283 1697
rect 1691 1657 3283 1663
rect -3339 1613 -3293 1625
rect -3339 637 -3333 1613
rect -3299 637 -3293 1613
rect -3339 625 -3293 637
rect -1681 1613 -1635 1625
rect -1681 637 -1675 1613
rect -1641 637 -1635 1613
rect -1681 625 -1635 637
rect -23 1613 23 1625
rect -23 637 -17 1613
rect 17 637 23 1613
rect -23 625 23 637
rect 1635 1613 1681 1625
rect 1635 637 1641 1613
rect 1675 637 1681 1613
rect 1635 625 1681 637
rect 3293 1613 3339 1625
rect 3293 637 3299 1613
rect 3333 637 3339 1613
rect 3293 625 3339 637
rect -3283 541 -1691 547
rect -3283 507 -3271 541
rect -1703 507 -1691 541
rect -3283 501 -1691 507
rect -1625 541 -33 547
rect -1625 507 -1613 541
rect -45 507 -33 541
rect -1625 501 -33 507
rect 33 541 1625 547
rect 33 507 45 541
rect 1613 507 1625 541
rect 33 501 1625 507
rect 1691 541 3283 547
rect 1691 507 1703 541
rect 3271 507 3283 541
rect 1691 501 3283 507
rect -3339 457 -3293 469
rect -3339 -519 -3333 457
rect -3299 -519 -3293 457
rect -3339 -531 -3293 -519
rect -1681 457 -1635 469
rect -1681 -519 -1675 457
rect -1641 -519 -1635 457
rect -1681 -531 -1635 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 1635 457 1681 469
rect 1635 -519 1641 457
rect 1675 -519 1681 457
rect 1635 -531 1681 -519
rect 3293 457 3339 469
rect 3293 -519 3299 457
rect 3333 -519 3339 457
rect 3293 -531 3339 -519
rect -3283 -615 -1691 -609
rect -3283 -649 -3271 -615
rect -1703 -649 -1691 -615
rect -3283 -655 -1691 -649
rect -1625 -615 -33 -609
rect -1625 -649 -1613 -615
rect -45 -649 -33 -615
rect -1625 -655 -33 -649
rect 33 -615 1625 -609
rect 33 -649 45 -615
rect 1613 -649 1625 -615
rect 33 -655 1625 -649
rect 1691 -615 3283 -609
rect 1691 -649 1703 -615
rect 3271 -649 3283 -615
rect 1691 -655 3283 -649
rect -3339 -699 -3293 -687
rect -3339 -1675 -3333 -699
rect -3299 -1675 -3293 -699
rect -3339 -1687 -3293 -1675
rect -1681 -699 -1635 -687
rect -1681 -1675 -1675 -699
rect -1641 -1675 -1635 -699
rect -1681 -1687 -1635 -1675
rect -23 -699 23 -687
rect -23 -1675 -17 -699
rect 17 -1675 23 -699
rect -23 -1687 23 -1675
rect 1635 -699 1681 -687
rect 1635 -1675 1641 -699
rect 1675 -1675 1681 -699
rect 1635 -1687 1681 -1675
rect 3293 -699 3339 -687
rect 3293 -1675 3299 -699
rect 3333 -1675 3339 -699
rect 3293 -1687 3339 -1675
rect -3283 -1771 -1691 -1765
rect -3283 -1805 -3271 -1771
rect -1703 -1805 -1691 -1771
rect -3283 -1811 -1691 -1805
rect -1625 -1771 -33 -1765
rect -1625 -1805 -1613 -1771
rect -45 -1805 -33 -1771
rect -1625 -1811 -33 -1805
rect 33 -1771 1625 -1765
rect 33 -1805 45 -1771
rect 1613 -1805 1625 -1771
rect 33 -1811 1625 -1805
rect 1691 -1771 3283 -1765
rect 1691 -1805 1703 -1771
rect 3271 -1805 3283 -1771
rect 1691 -1811 3283 -1805
rect -3339 -1855 -3293 -1843
rect -3339 -2831 -3333 -1855
rect -3299 -2831 -3293 -1855
rect -3339 -2843 -3293 -2831
rect -1681 -1855 -1635 -1843
rect -1681 -2831 -1675 -1855
rect -1641 -2831 -1635 -1855
rect -1681 -2843 -1635 -2831
rect -23 -1855 23 -1843
rect -23 -2831 -17 -1855
rect 17 -2831 23 -1855
rect -23 -2843 23 -2831
rect 1635 -1855 1681 -1843
rect 1635 -2831 1641 -1855
rect 1675 -2831 1681 -1855
rect 1635 -2843 1681 -2831
rect 3293 -1855 3339 -1843
rect 3293 -2831 3299 -1855
rect 3333 -2831 3339 -1855
rect 3293 -2843 3339 -2831
<< properties >>
string FIXED_BBOX -3450 -2974 3450 2974
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 8 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
