magic
tech sky130A
magscale 1 2
timestamp 1711689217
<< dnwell >>
rect -6407 -5578 10340 5402
<< nwell >>
rect -6487 5196 10420 5482
rect -6487 -5372 -6201 5196
rect 10134 -5372 10420 5196
rect -6487 -5658 10420 -5372
<< nsubdiff >>
rect -6450 5425 10383 5445
rect -6450 5391 -6370 5425
rect 10303 5391 10383 5425
rect -6450 5371 10383 5391
rect -6450 5365 -6376 5371
rect -6450 -5541 -6430 5365
rect -6396 -5541 -6376 5365
rect -6450 -5547 -6376 -5541
rect 10309 5365 10383 5371
rect 10309 -5541 10329 5365
rect 10363 -5541 10383 5365
rect 10309 -5547 10383 -5541
rect -6450 -5567 10383 -5547
rect -6450 -5601 -6370 -5567
rect 10303 -5601 10383 -5567
rect -6450 -5621 10383 -5601
<< nsubdiffcont >>
rect -6370 5391 10303 5425
rect -6430 -5541 -6396 5365
rect 10329 -5541 10363 5365
rect -6370 -5601 10303 -5567
<< locali >>
rect -67 6626 36 6671
rect -6430 5391 -6370 5425
rect 10303 5391 10363 5425
rect -6430 5365 -6396 5391
rect 10329 5365 10363 5391
rect -6430 -5567 -6396 -5541
rect 10329 -5567 10363 -5541
rect -6430 -5601 10363 -5567
<< viali >>
rect 100 -53 134 -19
rect 3416 -53 3450 -19
<< metal1 >>
rect -347 6493 -343 6539
rect -399 6461 -353 6465
rect -241 6461 -195 6465
rect 1742 451 1808 497
rect 91 407 143 419
rect 91 335 143 347
rect 1749 407 1801 419
rect 1749 335 1801 347
rect 3407 407 3459 419
rect 3407 335 3459 347
rect 1742 211 1808 257
rect 91 167 143 179
rect 91 95 143 107
rect 1749 167 1801 179
rect 1749 95 1801 107
rect 3407 167 3459 179
rect 3407 95 3459 107
rect 85 -6 149 0
rect 85 -66 91 -6
rect 143 -66 149 -6
rect 85 -72 149 -66
rect 3401 -6 3465 0
rect 3401 -66 3407 -6
rect 3459 -66 3465 -6
rect 3401 -72 3465 -66
<< via1 >>
rect 91 347 143 407
rect 1749 347 1801 407
rect 3407 347 3459 407
rect 91 107 143 167
rect 1749 107 1801 167
rect 3407 107 3459 167
rect 91 -19 143 -6
rect 91 -53 100 -19
rect 100 -53 134 -19
rect 134 -53 143 -19
rect 91 -66 143 -53
rect 3407 -19 3459 -6
rect 3407 -53 3416 -19
rect 3416 -53 3450 -19
rect 3450 -53 3459 -19
rect 3407 -66 3459 -53
<< metal2 >>
rect 91 407 143 419
rect 91 167 143 347
rect 1749 407 1801 419
rect 1749 335 1801 347
rect 3407 407 3459 419
rect 91 -6 143 107
rect 1749 167 1801 179
rect 1749 95 1801 107
rect 3407 167 3459 347
rect 91 -82 143 -66
rect 3407 -6 3459 107
rect 3407 -82 3459 -66
use sky130_fd_pr__nfet_g5v0d10v5_DHXKC7  sky130_fd_pr__nfet_g5v0d10v5_DHXKC7_0
timestamp 1711689129
transform 1 0 -297 0 1 6419
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_H4GRF3  sky130_fd_pr__nfet_g5v0d10v5_H4GRF3_0
timestamp 1711687497
transform 1 0 1775 0 1 288
box -1857 -389 1857 389
<< labels >>
rlabel metal1 1749 451 1749 451 5 vinn
rlabel metal2 1749 419 1749 419 1 vnn
rlabel metal2 1749 179 1749 179 1 vpp
rlabel metal1 1749 211 1749 211 5 vinp
rlabel metal2 91 279 91 279 7 vt
rlabel locali -6430 -5601 -6430 -5601 7 avdd
rlabel locali 36 6671 36 6671 1 avss
rlabel metal1 -399 6461 -399 6461 1 dd
rlabel metal1 -241 6461 -241 6461 1 ss
rlabel metal1 -343 6539 -343 6539 1 gg
<< end >>
