magic
tech sky130A
magscale 1 2
timestamp 1711687497
<< pwell >>
rect -1857 -389 1857 389
<< mvnmos >>
rect -1629 47 -29 131
rect 29 47 1629 131
rect -1629 -193 -29 -109
rect 29 -193 1629 -109
<< mvndiff >>
rect -1687 119 -1629 131
rect -1687 59 -1675 119
rect -1641 59 -1629 119
rect -1687 47 -1629 59
rect -29 119 29 131
rect -29 59 -17 119
rect 17 59 29 119
rect -29 47 29 59
rect 1629 119 1687 131
rect 1629 59 1641 119
rect 1675 59 1687 119
rect 1629 47 1687 59
rect -1687 -121 -1629 -109
rect -1687 -181 -1675 -121
rect -1641 -181 -1629 -121
rect -1687 -193 -1629 -181
rect -29 -121 29 -109
rect -29 -181 -17 -121
rect 17 -181 29 -121
rect -29 -193 29 -181
rect 1629 -121 1687 -109
rect 1629 -181 1641 -121
rect 1675 -181 1687 -121
rect 1629 -193 1687 -181
<< mvndiffc >>
rect -1675 59 -1641 119
rect -17 59 17 119
rect 1641 59 1675 119
rect -1675 -181 -1641 -121
rect -17 -181 17 -121
rect 1641 -181 1675 -121
<< mvpsubdiff >>
rect -1821 341 1821 353
rect -1821 307 -1713 341
rect 1713 307 1821 341
rect -1821 295 1821 307
rect -1821 245 -1763 295
rect -1821 -245 -1809 245
rect -1775 -245 -1763 245
rect 1763 245 1821 295
rect -1821 -295 -1763 -245
rect 1763 -245 1775 245
rect 1809 -245 1821 245
rect 1763 -295 1821 -245
rect -1821 -307 1821 -295
rect -1821 -341 -1713 -307
rect 1713 -341 1821 -307
rect -1821 -353 1821 -341
<< mvpsubdiffcont >>
rect -1713 307 1713 341
rect -1809 -245 -1775 245
rect 1775 -245 1809 245
rect -1713 -341 1713 -307
<< poly >>
rect -1629 203 -29 219
rect -1629 169 -1613 203
rect -45 169 -29 203
rect -1629 131 -29 169
rect 29 203 1629 219
rect 29 169 45 203
rect 1613 169 1629 203
rect 29 131 1629 169
rect -1629 21 -29 47
rect 29 21 1629 47
rect -1629 -37 -29 -21
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect -1629 -109 -29 -71
rect 29 -37 1629 -21
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect 29 -109 1629 -71
rect -1629 -219 -29 -193
rect 29 -219 1629 -193
<< polycont >>
rect -1613 169 -45 203
rect 45 169 1613 203
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
<< locali >>
rect -1809 307 -1713 341
rect 1713 307 1809 341
rect -1809 245 -1775 307
rect 1775 245 1809 307
rect -1629 169 -1613 203
rect -45 169 -29 203
rect 29 169 45 203
rect 1613 169 1629 203
rect -1675 119 -1641 135
rect -1675 43 -1641 59
rect -17 119 17 135
rect -17 43 17 59
rect 1641 119 1675 135
rect 1641 43 1675 59
rect -1629 -71 -1613 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1613 -71 1629 -37
rect -1675 -121 -1641 -105
rect -1675 -197 -1641 -181
rect -17 -121 17 -105
rect -17 -197 17 -181
rect 1641 -121 1675 -105
rect 1641 -197 1675 -181
rect -1809 -307 -1775 -245
rect 1775 -307 1809 -245
rect -1809 -341 -1713 -307
rect 1713 -341 1809 -307
<< viali >>
rect -1613 169 -45 203
rect 45 169 1613 203
rect -1675 59 -1641 119
rect -17 59 17 119
rect 1641 59 1675 119
rect -1613 -71 -45 -37
rect 45 -71 1613 -37
rect -1675 -181 -1641 -121
rect -17 -181 17 -121
rect 1641 -181 1675 -121
<< metal1 >>
rect -1625 203 -33 209
rect -1625 169 -1613 203
rect -45 169 -33 203
rect -1625 163 -33 169
rect 33 203 1625 209
rect 33 169 45 203
rect 1613 169 1625 203
rect 33 163 1625 169
rect -1681 119 -1635 131
rect -1681 59 -1675 119
rect -1641 59 -1635 119
rect -1681 47 -1635 59
rect -23 119 23 131
rect -23 59 -17 119
rect 17 59 23 119
rect -23 47 23 59
rect 1635 119 1681 131
rect 1635 59 1641 119
rect 1675 59 1681 119
rect 1635 47 1681 59
rect -1625 -37 -33 -31
rect -1625 -71 -1613 -37
rect -45 -71 -33 -37
rect -1625 -77 -33 -71
rect 33 -37 1625 -31
rect 33 -71 45 -37
rect 1613 -71 1625 -37
rect 33 -77 1625 -71
rect -1681 -121 -1635 -109
rect -1681 -181 -1675 -121
rect -1641 -181 -1635 -121
rect -1681 -193 -1635 -181
rect -23 -121 23 -109
rect -23 -181 -17 -121
rect 17 -181 23 -121
rect -23 -193 23 -181
rect 1635 -121 1681 -109
rect 1635 -181 1641 -121
rect 1675 -181 1681 -121
rect 1635 -193 1681 -181
<< properties >>
string FIXED_BBOX -1792 -324 1792 324
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 8 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
