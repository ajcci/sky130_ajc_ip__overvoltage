magic
tech sky130A
magscale 1 2
timestamp 1712165136
<< error_s >>
rect 10441 7207 10515 7216
rect 10441 7151 10450 7207
rect 10441 7142 10515 7151
rect 9958 6959 10032 6968
rect 10441 6959 10515 6968
rect 9958 6903 9967 6959
rect 10441 6903 10450 6959
rect 9958 6894 10032 6903
rect 10441 6894 10515 6903
<< locali >>
rect 12546 8650 12610 8665
rect 12546 8616 12561 8650
rect 12595 8616 12610 8650
rect 12546 8601 12610 8616
rect 12701 8644 12765 8659
rect 12701 8546 12716 8644
rect 12750 8546 12765 8644
rect 12701 8531 12765 8546
rect 12965 7927 13085 8032
rect 10237 7265 10365 7280
rect 10237 7167 10252 7265
rect 10350 7167 10365 7265
rect 10581 7265 10645 7280
rect 10237 7152 10365 7167
rect 10446 7196 10510 7211
rect 10446 7162 10461 7196
rect 10495 7162 10510 7196
rect 10446 7147 10510 7162
rect 10581 7167 10596 7265
rect 10630 7167 10645 7265
rect 10581 7152 10645 7167
rect 11317 7149 11375 7161
rect 11317 7115 11329 7149
rect 11363 7115 11375 7149
rect 11317 7103 11375 7115
rect 11161 7007 11289 7022
rect 11161 6909 11176 7007
rect 11274 6909 11289 7007
rect 11429 7007 11493 7022
rect 11161 6894 11289 6909
rect 11330 6943 11394 6958
rect 11330 6909 11345 6943
rect 11379 6909 11394 6943
rect 11330 6894 11394 6909
rect 11429 6909 11444 7007
rect 11478 6909 11493 7007
rect 11429 6894 11493 6909
rect 11275 6639 11403 6654
rect 11275 6605 11290 6639
rect 11388 6605 11403 6639
rect 11275 6590 11403 6605
<< viali >>
rect 12561 8616 12595 8650
rect 12716 8546 12750 8644
rect 10252 7167 10350 7265
rect 10461 7162 10495 7196
rect 10596 7167 10630 7265
rect 11329 7115 11363 7149
rect 11176 6909 11274 7007
rect 11345 6909 11379 6943
rect 11444 6909 11478 7007
rect 11290 6605 11388 6639
<< metal1 >>
rect 12546 8659 12610 8665
rect 12546 8607 12552 8659
rect 12604 8607 12610 8659
rect 12546 8601 12610 8607
rect 12701 8653 12765 8659
rect 12701 8537 12707 8653
rect 12759 8537 12765 8653
rect 12701 8531 12765 8537
rect 12661 7945 12725 7951
rect 12661 7893 12667 7945
rect 12719 7933 12725 7945
rect 12719 7893 12791 7933
rect 12661 7887 12791 7893
rect 10227 7279 10375 7290
rect 10227 7153 10238 7279
rect 10364 7153 10375 7279
rect 10576 7279 10650 7290
rect 10227 7142 10375 7153
rect 10441 7205 10515 7216
rect 10441 7153 10452 7205
rect 10504 7153 10515 7205
rect 10441 7142 10515 7153
rect 10576 7153 10587 7279
rect 10639 7153 10650 7279
rect 10576 7142 10650 7153
rect 11317 7149 11375 7161
rect 11317 7115 11329 7149
rect 11363 7115 11375 7149
rect 11317 7103 11375 7115
rect 12640 7098 12704 7102
rect 12602 7096 12704 7098
rect 12602 7044 12646 7096
rect 12698 7044 12704 7096
rect 12602 7042 12704 7044
rect 10227 7031 10375 7042
rect 10227 6905 10238 7031
rect 10364 6905 10375 7031
rect 10576 7031 10650 7042
rect 12640 7038 12704 7042
rect 12904 7096 12968 7102
rect 10227 6894 10375 6905
rect 10441 6957 10515 6968
rect 10441 6905 10452 6957
rect 10504 6905 10515 6957
rect 10441 6894 10515 6905
rect 10576 6905 10587 7031
rect 10639 6905 10650 7031
rect 10576 6894 10650 6905
rect 10733 7016 10861 7022
rect 10733 6900 10739 7016
rect 10855 6900 10861 7016
rect 11001 7016 11065 7022
rect 10733 6894 10861 6900
rect 10902 6952 10966 6958
rect 10902 6900 10908 6952
rect 10960 6900 10966 6952
rect 10902 6894 10966 6900
rect 11001 6900 11007 7016
rect 11059 6900 11065 7016
rect 11001 6894 11065 6900
rect 11161 7016 11289 7022
rect 11161 6900 11167 7016
rect 11283 6900 11289 7016
rect 11429 7016 11493 7022
rect 11161 6894 11289 6900
rect 11330 6952 11394 6958
rect 11330 6900 11336 6952
rect 11388 6900 11394 6952
rect 11330 6894 11394 6900
rect 11429 6900 11435 7016
rect 11487 6900 11493 7016
rect 12904 6980 12910 7096
rect 12962 6980 12968 7096
rect 12904 6974 12968 6980
rect 11429 6894 11493 6900
rect 12726 6968 12790 6974
rect 12726 6852 12732 6968
rect 12784 6852 12790 6968
rect 12726 6846 12790 6852
rect 11021 6722 11149 6728
rect 11021 6670 11027 6722
rect 11143 6670 11149 6722
rect 11021 6664 11149 6670
rect 11275 6648 11403 6654
rect 10585 6633 10733 6644
rect 10585 6581 10596 6633
rect 10722 6581 10733 6633
rect 11275 6596 11281 6648
rect 11397 6596 11403 6648
rect 11275 6590 11403 6596
rect 10585 6570 10733 6581
rect 12548 6385 12676 6391
rect 12548 6333 12554 6385
rect 12670 6333 12676 6385
rect 12548 6327 12676 6333
rect 12725 6327 12791 6373
rect 12726 6289 12790 6295
rect 12548 6182 12612 6188
rect 12548 6066 12554 6182
rect 12606 6066 12612 6182
rect 12726 6173 12732 6289
rect 12784 6173 12790 6289
rect 12726 6167 12790 6173
rect 12904 6182 12968 6188
rect 12548 6060 12612 6066
rect 12904 6066 12910 6182
rect 12962 6066 12968 6182
rect 12904 6060 12968 6066
rect 784 4059 900 4480
rect 1540 4059 1656 4480
rect 2296 4059 2412 4480
rect 3052 4059 3168 4480
rect 3808 4059 3924 4480
rect 4564 4059 4680 4480
rect 5320 4059 5436 4480
rect 6076 4059 6192 4480
rect 6832 4059 6948 4480
rect 7588 4059 7704 4480
rect 8344 4059 8460 4480
rect 9100 4059 9216 4480
rect 9856 4059 9972 4480
rect 10612 4059 10728 4480
rect 11368 4059 11484 4480
rect 12124 4059 12240 4480
rect 12880 4059 12996 4480
rect 13636 4059 13752 4480
rect 14392 4059 14508 4480
rect 15148 4059 15264 4480
rect 15904 4059 16020 4480
rect 16660 4059 16776 4480
rect 17416 4059 17532 4480
rect 18172 4059 18288 4480
rect 18928 4059 19044 4480
rect 19684 4059 19800 4480
rect 20440 4059 20556 4480
rect 21196 4059 21312 4480
rect 21952 4059 22068 4480
rect 22708 4059 22824 4480
rect 23464 4059 23580 4480
rect 24220 4059 24336 4480
rect 24976 4059 25092 4480
rect 25732 4059 25848 4480
rect 26488 4059 26604 4480
rect 27244 4059 27360 4480
rect 28000 4059 28116 4480
rect 28756 4059 28872 4480
rect 29512 4059 29628 4480
rect 30268 4059 30384 4480
rect 31024 4059 31140 4480
rect 31780 4059 31896 4480
rect 32536 4059 32652 4480
rect 33292 4059 33408 4480
rect 34048 4059 34164 4480
rect 34804 4059 34920 4480
rect 35560 4059 35676 4480
rect 36316 4059 36432 4480
rect 37072 4059 37188 4480
rect 37828 4059 37944 4480
rect 38584 4059 38700 4480
rect 39340 4059 39456 4480
rect 406 140 522 561
rect 1162 140 1278 561
rect 1918 140 2034 561
rect 2674 140 2790 561
rect 3430 140 3546 561
rect 4186 140 4302 561
rect 4942 140 5058 561
rect 5698 140 5814 561
rect 6454 140 6570 561
rect 7210 140 7326 561
rect 7966 140 8082 561
rect 8722 140 8838 561
rect 9478 140 9594 561
rect 10234 140 10350 561
rect 10990 140 11106 561
rect 11746 140 11862 561
rect 12502 140 12618 561
rect 13258 140 13374 561
rect 14014 140 14130 561
rect 14770 140 14886 561
rect 15526 140 15642 561
rect 16282 140 16398 561
rect 17038 140 17154 561
rect 17794 140 17910 561
rect 18550 140 18666 561
rect 19306 140 19422 561
rect 20062 140 20178 561
rect 20818 140 20934 561
rect 21574 140 21690 561
rect 22330 140 22446 561
rect 23086 140 23202 561
rect 23842 140 23958 561
rect 24598 140 24714 561
rect 25354 140 25470 561
rect 26110 140 26226 561
rect 26866 140 26982 561
rect 27622 140 27738 561
rect 28378 140 28494 561
rect 29134 140 29250 561
rect 29890 140 30006 561
rect 30646 140 30762 561
rect 31402 140 31518 561
rect 32158 140 32274 561
rect 32914 140 33030 561
rect 33670 140 33786 561
rect 34426 140 34542 561
rect 35182 140 35298 561
rect 35938 140 36054 561
rect 36694 140 36810 561
rect 37450 140 37566 561
rect 38206 140 38322 561
rect 38962 140 39078 561
<< via1 >>
rect 12552 8650 12604 8659
rect 12552 8616 12561 8650
rect 12561 8616 12595 8650
rect 12595 8616 12604 8650
rect 12552 8607 12604 8616
rect 12707 8644 12759 8653
rect 12707 8546 12716 8644
rect 12716 8546 12750 8644
rect 12750 8546 12759 8644
rect 12707 8537 12759 8546
rect 12667 7893 12719 7945
rect 10238 7265 10364 7279
rect 10238 7167 10252 7265
rect 10252 7167 10350 7265
rect 10350 7167 10364 7265
rect 10238 7153 10364 7167
rect 10452 7196 10504 7205
rect 10452 7162 10461 7196
rect 10461 7162 10495 7196
rect 10495 7162 10504 7196
rect 10452 7153 10504 7162
rect 10587 7265 10639 7279
rect 10587 7167 10596 7265
rect 10596 7167 10630 7265
rect 10630 7167 10639 7265
rect 10587 7153 10639 7167
rect 12646 7044 12698 7096
rect 10238 6905 10364 7031
rect 10452 6905 10504 6957
rect 10587 6905 10639 7031
rect 10739 6900 10855 7016
rect 10908 6900 10960 6952
rect 11007 6900 11059 7016
rect 11167 7007 11283 7016
rect 11167 6909 11176 7007
rect 11176 6909 11274 7007
rect 11274 6909 11283 7007
rect 11167 6900 11283 6909
rect 11336 6943 11388 6952
rect 11336 6909 11345 6943
rect 11345 6909 11379 6943
rect 11379 6909 11388 6943
rect 11336 6900 11388 6909
rect 11435 7007 11487 7016
rect 11435 6909 11444 7007
rect 11444 6909 11478 7007
rect 11478 6909 11487 7007
rect 11435 6900 11487 6909
rect 12910 6980 12962 7096
rect 12732 6852 12784 6968
rect 11027 6670 11143 6722
rect 10596 6581 10722 6633
rect 11281 6639 11397 6648
rect 11281 6605 11290 6639
rect 11290 6605 11388 6639
rect 11388 6605 11397 6639
rect 11281 6596 11397 6605
rect 12554 6333 12670 6385
rect 12554 6066 12606 6182
rect 12732 6173 12784 6289
rect 12910 6066 12962 6182
<< metal2 >>
rect 12546 8659 12610 8665
rect 12546 8607 12552 8659
rect 12604 8607 12610 8659
rect 12546 8601 12610 8607
rect 12701 8653 12765 8659
rect 10227 7281 10375 7290
rect 10227 7151 10236 7281
rect 10366 7151 10375 7281
rect 10576 7281 10650 7290
rect 10227 7142 10375 7151
rect 10441 7207 10515 7216
rect 10441 7151 10450 7207
rect 10506 7151 10515 7207
rect 10441 7142 10515 7151
rect 10576 7151 10585 7281
rect 10641 7151 10650 7281
rect 10576 7142 10650 7151
rect 9743 7033 9891 7042
rect 9743 6903 9752 7033
rect 9882 6903 9891 7033
rect 10092 7033 10166 7042
rect 9743 6894 9891 6903
rect 9958 6959 10032 6968
rect 9958 6903 9967 6959
rect 10023 6903 10032 6959
rect 9958 6894 10032 6903
rect 10092 6903 10101 7033
rect 10157 6903 10166 7033
rect 10092 6894 10166 6903
rect 10227 7033 10375 7042
rect 10227 6903 10236 7033
rect 10366 6903 10375 7033
rect 10576 7033 10650 7042
rect 10227 6894 10375 6903
rect 10441 6959 10515 6968
rect 10441 6903 10450 6959
rect 10506 6903 10515 6959
rect 10441 6894 10515 6903
rect 10576 6903 10585 7033
rect 10641 6903 10650 7033
rect 10576 6894 10650 6903
rect 10733 7016 10861 7022
rect 10733 6900 10739 7016
rect 10855 6900 10861 7016
rect 11001 7016 11065 7022
rect 10733 6894 10861 6900
rect 10902 6952 10966 6958
rect 10902 6900 10908 6952
rect 10960 6900 10966 6952
rect 10902 6894 10966 6900
rect 11001 6900 11007 7016
rect 11059 6900 11065 7016
rect 11001 6894 11065 6900
rect 11161 7016 11289 7022
rect 11161 6900 11167 7016
rect 11283 6900 11289 7016
rect 11429 7016 11493 7022
rect 11161 6894 11289 6900
rect 11330 6952 11394 6958
rect 11330 6900 11336 6952
rect 11388 6900 11394 6952
rect 11330 6894 11394 6900
rect 11429 6900 11435 7016
rect 11487 6900 11493 7016
rect 11429 6894 11493 6900
rect 11021 6722 11149 6728
rect 10101 6679 10249 6688
rect 10101 6623 10110 6679
rect 10240 6623 10249 6679
rect 11021 6670 11027 6722
rect 11143 6670 11149 6722
rect 11021 6664 11149 6670
rect 11275 6648 11403 6654
rect 10101 6614 10249 6623
rect 10585 6635 10733 6644
rect 10585 6579 10594 6635
rect 10724 6579 10733 6635
rect 11275 6596 11281 6648
rect 11397 6596 11403 6648
rect 11275 6590 11403 6596
rect 10585 6570 10733 6579
rect 12552 6391 12608 8601
rect 12701 8581 12707 8653
rect 12664 8537 12707 8581
rect 12759 8537 12765 8653
rect 12664 8531 12765 8537
rect 12664 7951 12720 8531
rect 12661 7945 12725 7951
rect 12661 7893 12667 7945
rect 12719 7893 12725 7945
rect 12661 7887 12725 7893
rect 12640 7098 12704 7102
rect 12904 7098 12968 7102
rect 12640 7096 12968 7098
rect 12640 7044 12646 7096
rect 12698 7044 12910 7096
rect 12640 7042 12910 7044
rect 12640 7038 12704 7042
rect 12904 6980 12910 7042
rect 12962 6980 12968 7096
rect 12904 6974 12968 6980
rect 12726 6968 12790 6974
rect 12726 6852 12732 6968
rect 12784 6852 12790 6968
rect 12726 6846 12790 6852
rect 12548 6385 12676 6391
rect 12548 6333 12554 6385
rect 12670 6333 12676 6385
rect 12548 6327 12676 6333
rect 12730 6295 12786 6846
rect 12726 6289 12790 6295
rect 12548 6182 12612 6188
rect 12548 6066 12554 6182
rect 12606 6116 12612 6182
rect 12726 6173 12732 6289
rect 12784 6173 12790 6289
rect 12908 6188 12964 6974
rect 12726 6167 12790 6173
rect 12904 6182 12968 6188
rect 12904 6116 12910 6182
rect 12606 6066 12910 6116
rect 12962 6066 12968 6182
rect 12548 6060 12968 6066
<< via2 >>
rect 10236 7279 10366 7281
rect 10236 7153 10238 7279
rect 10238 7153 10364 7279
rect 10364 7153 10366 7279
rect 10236 7151 10366 7153
rect 10450 7205 10506 7207
rect 10450 7153 10452 7205
rect 10452 7153 10504 7205
rect 10504 7153 10506 7205
rect 10450 7151 10506 7153
rect 10585 7279 10641 7281
rect 10585 7153 10587 7279
rect 10587 7153 10639 7279
rect 10639 7153 10641 7279
rect 10585 7151 10641 7153
rect 9752 6903 9882 7033
rect 9967 6903 10023 6959
rect 10101 6903 10157 7033
rect 10236 7031 10366 7033
rect 10236 6905 10238 7031
rect 10238 6905 10364 7031
rect 10364 6905 10366 7031
rect 10236 6903 10366 6905
rect 10450 6957 10506 6959
rect 10450 6905 10452 6957
rect 10452 6905 10504 6957
rect 10504 6905 10506 6957
rect 10450 6903 10506 6905
rect 10585 7031 10641 7033
rect 10585 6905 10587 7031
rect 10587 6905 10639 7031
rect 10639 6905 10641 7031
rect 10585 6903 10641 6905
rect 10110 6623 10240 6679
rect 10594 6633 10724 6635
rect 10594 6581 10596 6633
rect 10596 6581 10722 6633
rect 10722 6581 10724 6633
rect 10594 6579 10724 6581
<< metal3 >>
rect 10227 7281 10375 7290
rect 10227 7151 10236 7281
rect 10366 7151 10375 7281
rect 10576 7281 10650 7290
rect 10227 7142 10375 7151
rect 10441 7207 10515 7216
rect 10441 7151 10450 7207
rect 10506 7151 10515 7207
rect 10441 7142 10515 7151
rect 10576 7151 10585 7281
rect 10641 7151 10650 7281
rect 10576 7142 10650 7151
rect 9743 7033 9891 7042
rect 9743 6903 9752 7033
rect 9882 6903 9891 7033
rect 10092 7033 10166 7042
rect 9743 6894 9891 6903
rect 9958 6959 10032 6968
rect 9958 6903 9967 6959
rect 10023 6903 10032 6959
rect 9958 6894 10032 6903
rect 10092 6903 10101 7033
rect 10157 6903 10166 7033
rect 10092 6894 10166 6903
rect 10227 7033 10375 7042
rect 10227 6903 10236 7033
rect 10366 6903 10375 7033
rect 10576 7033 10650 7042
rect 10227 6894 10375 6903
rect 10441 6959 10515 6968
rect 10441 6903 10450 6959
rect 10506 6903 10515 6959
rect 10441 6894 10515 6903
rect 10576 6903 10585 7033
rect 10641 6903 10650 7033
rect 10576 6894 10650 6903
rect 10101 6679 10249 6688
rect 10101 6623 10110 6679
rect 10240 6623 10249 6679
rect 10101 6614 10249 6623
rect 10585 6635 10733 6644
rect 10585 6579 10594 6635
rect 10724 6579 10733 6635
rect 10585 6570 10733 6579
use sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ  sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ_0
timestamp 1712160855
transform 1 0 16763 0 1 5826
box -4382 -727 4382 727
use sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY  sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY_0
timestamp 1712158818
transform 1 0 16763 0 1 7382
box -4412 -762 4412 762
use sky130_fd_pr__res_xhigh_po_1p41_CZUCEE  sky130_fd_pr__res_xhigh_po_1p41_CZUCEE_0
timestamp 1712156631
transform 1 0 19931 0 1 2310
box -19963 -2342 19963 2342
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1707688321
transform 1 0 12499 0 1 8285
box -66 -43 354 897
<< labels >>
flabel metal1 s 31034 4480 31034 4480 0 FreeSans 800 0 0 0 vtrip15
flabel metal1 s 30278 4480 30278 4480 0 FreeSans 800 0 0 0 vtrip13
flabel metal1 s 29522 4480 29522 4480 0 FreeSans 800 0 0 0 vtrip11
flabel metal1 s 28766 4480 28766 4480 0 FreeSans 800 0 0 0 vtrip9
flabel metal1 s 28010 4480 28010 4480 0 FreeSans 800 0 0 0 vtrip7
flabel metal1 s 27254 4480 27254 4480 0 FreeSans 800 0 0 0 vtrip5
flabel metal1 s 26498 4480 26498 4480 0 FreeSans 800 0 0 0 vtrip3
flabel metal1 s 25742 4480 25742 4480 0 FreeSans 800 0 0 0 vtrip1
flabel metal1 s 25364 140 25364 140 0 FreeSans 800 0 0 0 vtrip0
flabel metal1 s 26120 140 26120 140 0 FreeSans 800 0 0 0 vtrip2
flabel metal1 s 26876 140 26876 140 0 FreeSans 800 0 0 0 vtrip4
flabel metal1 s 27632 140 27632 140 0 FreeSans 800 0 0 0 vtrip6
flabel metal1 s 28388 140 28388 140 0 FreeSans 800 0 0 0 vtrip8
flabel metal1 s 29144 140 29144 140 0 FreeSans 800 0 0 0 vtrip10
flabel metal1 s 29900 140 29900 140 0 FreeSans 800 0 0 0 vtrip12
flabel metal1 s 30656 140 30656 140 0 FreeSans 800 0 0 0 vtrip14
<< end >>
