* SPICE3 file created from comparator_wip_flattened2.ext - technology: sky130A

.subckt comparator_wip_flattened2 avdd
X0 s g d vt sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
C0 avdd vt 1.02054p
C1 avdd avss 1.12261p
.ends
