magic
tech sky130A
magscale 1 2
timestamp 1712158818
<< nwell >>
rect -4412 -797 4412 797
<< mvpmos >>
rect -4154 -500 -4034 500
rect -3976 -500 -3856 500
rect -3798 -500 -3678 500
rect -3620 -500 -3500 500
rect -3442 -500 -3322 500
rect -3264 -500 -3144 500
rect -3086 -500 -2966 500
rect -2908 -500 -2788 500
rect -2730 -500 -2610 500
rect -2552 -500 -2432 500
rect -2374 -500 -2254 500
rect -2196 -500 -2076 500
rect -2018 -500 -1898 500
rect -1840 -500 -1720 500
rect -1662 -500 -1542 500
rect -1484 -500 -1364 500
rect -1306 -500 -1186 500
rect -1128 -500 -1008 500
rect -950 -500 -830 500
rect -772 -500 -652 500
rect -594 -500 -474 500
rect -416 -500 -296 500
rect -238 -500 -118 500
rect -60 -500 60 500
rect 118 -500 238 500
rect 296 -500 416 500
rect 474 -500 594 500
rect 652 -500 772 500
rect 830 -500 950 500
rect 1008 -500 1128 500
rect 1186 -500 1306 500
rect 1364 -500 1484 500
rect 1542 -500 1662 500
rect 1720 -500 1840 500
rect 1898 -500 2018 500
rect 2076 -500 2196 500
rect 2254 -500 2374 500
rect 2432 -500 2552 500
rect 2610 -500 2730 500
rect 2788 -500 2908 500
rect 2966 -500 3086 500
rect 3144 -500 3264 500
rect 3322 -500 3442 500
rect 3500 -500 3620 500
rect 3678 -500 3798 500
rect 3856 -500 3976 500
rect 4034 -500 4154 500
<< mvpdiff >>
rect -4212 488 -4154 500
rect -4212 -488 -4200 488
rect -4166 -488 -4154 488
rect -4212 -500 -4154 -488
rect -4034 488 -3976 500
rect -4034 -488 -4022 488
rect -3988 -488 -3976 488
rect -4034 -500 -3976 -488
rect -3856 488 -3798 500
rect -3856 -488 -3844 488
rect -3810 -488 -3798 488
rect -3856 -500 -3798 -488
rect -3678 488 -3620 500
rect -3678 -488 -3666 488
rect -3632 -488 -3620 488
rect -3678 -500 -3620 -488
rect -3500 488 -3442 500
rect -3500 -488 -3488 488
rect -3454 -488 -3442 488
rect -3500 -500 -3442 -488
rect -3322 488 -3264 500
rect -3322 -488 -3310 488
rect -3276 -488 -3264 488
rect -3322 -500 -3264 -488
rect -3144 488 -3086 500
rect -3144 -488 -3132 488
rect -3098 -488 -3086 488
rect -3144 -500 -3086 -488
rect -2966 488 -2908 500
rect -2966 -488 -2954 488
rect -2920 -488 -2908 488
rect -2966 -500 -2908 -488
rect -2788 488 -2730 500
rect -2788 -488 -2776 488
rect -2742 -488 -2730 488
rect -2788 -500 -2730 -488
rect -2610 488 -2552 500
rect -2610 -488 -2598 488
rect -2564 -488 -2552 488
rect -2610 -500 -2552 -488
rect -2432 488 -2374 500
rect -2432 -488 -2420 488
rect -2386 -488 -2374 488
rect -2432 -500 -2374 -488
rect -2254 488 -2196 500
rect -2254 -488 -2242 488
rect -2208 -488 -2196 488
rect -2254 -500 -2196 -488
rect -2076 488 -2018 500
rect -2076 -488 -2064 488
rect -2030 -488 -2018 488
rect -2076 -500 -2018 -488
rect -1898 488 -1840 500
rect -1898 -488 -1886 488
rect -1852 -488 -1840 488
rect -1898 -500 -1840 -488
rect -1720 488 -1662 500
rect -1720 -488 -1708 488
rect -1674 -488 -1662 488
rect -1720 -500 -1662 -488
rect -1542 488 -1484 500
rect -1542 -488 -1530 488
rect -1496 -488 -1484 488
rect -1542 -500 -1484 -488
rect -1364 488 -1306 500
rect -1364 -488 -1352 488
rect -1318 -488 -1306 488
rect -1364 -500 -1306 -488
rect -1186 488 -1128 500
rect -1186 -488 -1174 488
rect -1140 -488 -1128 488
rect -1186 -500 -1128 -488
rect -1008 488 -950 500
rect -1008 -488 -996 488
rect -962 -488 -950 488
rect -1008 -500 -950 -488
rect -830 488 -772 500
rect -830 -488 -818 488
rect -784 -488 -772 488
rect -830 -500 -772 -488
rect -652 488 -594 500
rect -652 -488 -640 488
rect -606 -488 -594 488
rect -652 -500 -594 -488
rect -474 488 -416 500
rect -474 -488 -462 488
rect -428 -488 -416 488
rect -474 -500 -416 -488
rect -296 488 -238 500
rect -296 -488 -284 488
rect -250 -488 -238 488
rect -296 -500 -238 -488
rect -118 488 -60 500
rect -118 -488 -106 488
rect -72 -488 -60 488
rect -118 -500 -60 -488
rect 60 488 118 500
rect 60 -488 72 488
rect 106 -488 118 488
rect 60 -500 118 -488
rect 238 488 296 500
rect 238 -488 250 488
rect 284 -488 296 488
rect 238 -500 296 -488
rect 416 488 474 500
rect 416 -488 428 488
rect 462 -488 474 488
rect 416 -500 474 -488
rect 594 488 652 500
rect 594 -488 606 488
rect 640 -488 652 488
rect 594 -500 652 -488
rect 772 488 830 500
rect 772 -488 784 488
rect 818 -488 830 488
rect 772 -500 830 -488
rect 950 488 1008 500
rect 950 -488 962 488
rect 996 -488 1008 488
rect 950 -500 1008 -488
rect 1128 488 1186 500
rect 1128 -488 1140 488
rect 1174 -488 1186 488
rect 1128 -500 1186 -488
rect 1306 488 1364 500
rect 1306 -488 1318 488
rect 1352 -488 1364 488
rect 1306 -500 1364 -488
rect 1484 488 1542 500
rect 1484 -488 1496 488
rect 1530 -488 1542 488
rect 1484 -500 1542 -488
rect 1662 488 1720 500
rect 1662 -488 1674 488
rect 1708 -488 1720 488
rect 1662 -500 1720 -488
rect 1840 488 1898 500
rect 1840 -488 1852 488
rect 1886 -488 1898 488
rect 1840 -500 1898 -488
rect 2018 488 2076 500
rect 2018 -488 2030 488
rect 2064 -488 2076 488
rect 2018 -500 2076 -488
rect 2196 488 2254 500
rect 2196 -488 2208 488
rect 2242 -488 2254 488
rect 2196 -500 2254 -488
rect 2374 488 2432 500
rect 2374 -488 2386 488
rect 2420 -488 2432 488
rect 2374 -500 2432 -488
rect 2552 488 2610 500
rect 2552 -488 2564 488
rect 2598 -488 2610 488
rect 2552 -500 2610 -488
rect 2730 488 2788 500
rect 2730 -488 2742 488
rect 2776 -488 2788 488
rect 2730 -500 2788 -488
rect 2908 488 2966 500
rect 2908 -488 2920 488
rect 2954 -488 2966 488
rect 2908 -500 2966 -488
rect 3086 488 3144 500
rect 3086 -488 3098 488
rect 3132 -488 3144 488
rect 3086 -500 3144 -488
rect 3264 488 3322 500
rect 3264 -488 3276 488
rect 3310 -488 3322 488
rect 3264 -500 3322 -488
rect 3442 488 3500 500
rect 3442 -488 3454 488
rect 3488 -488 3500 488
rect 3442 -500 3500 -488
rect 3620 488 3678 500
rect 3620 -488 3632 488
rect 3666 -488 3678 488
rect 3620 -500 3678 -488
rect 3798 488 3856 500
rect 3798 -488 3810 488
rect 3844 -488 3856 488
rect 3798 -500 3856 -488
rect 3976 488 4034 500
rect 3976 -488 3988 488
rect 4022 -488 4034 488
rect 3976 -500 4034 -488
rect 4154 488 4212 500
rect 4154 -488 4166 488
rect 4200 -488 4212 488
rect 4154 -500 4212 -488
<< mvpdiffc >>
rect -4200 -488 -4166 488
rect -4022 -488 -3988 488
rect -3844 -488 -3810 488
rect -3666 -488 -3632 488
rect -3488 -488 -3454 488
rect -3310 -488 -3276 488
rect -3132 -488 -3098 488
rect -2954 -488 -2920 488
rect -2776 -488 -2742 488
rect -2598 -488 -2564 488
rect -2420 -488 -2386 488
rect -2242 -488 -2208 488
rect -2064 -488 -2030 488
rect -1886 -488 -1852 488
rect -1708 -488 -1674 488
rect -1530 -488 -1496 488
rect -1352 -488 -1318 488
rect -1174 -488 -1140 488
rect -996 -488 -962 488
rect -818 -488 -784 488
rect -640 -488 -606 488
rect -462 -488 -428 488
rect -284 -488 -250 488
rect -106 -488 -72 488
rect 72 -488 106 488
rect 250 -488 284 488
rect 428 -488 462 488
rect 606 -488 640 488
rect 784 -488 818 488
rect 962 -488 996 488
rect 1140 -488 1174 488
rect 1318 -488 1352 488
rect 1496 -488 1530 488
rect 1674 -488 1708 488
rect 1852 -488 1886 488
rect 2030 -488 2064 488
rect 2208 -488 2242 488
rect 2386 -488 2420 488
rect 2564 -488 2598 488
rect 2742 -488 2776 488
rect 2920 -488 2954 488
rect 3098 -488 3132 488
rect 3276 -488 3310 488
rect 3454 -488 3488 488
rect 3632 -488 3666 488
rect 3810 -488 3844 488
rect 3988 -488 4022 488
rect 4166 -488 4200 488
<< mvnsubdiff >>
rect -4346 719 4346 731
rect -4346 685 -4238 719
rect 4238 685 4346 719
rect -4346 673 4346 685
rect -4346 623 -4288 673
rect -4346 -623 -4334 623
rect -4300 -623 -4288 623
rect 4288 623 4346 673
rect -4346 -673 -4288 -623
rect 4288 -623 4300 623
rect 4334 -623 4346 623
rect 4288 -673 4346 -623
rect -4346 -685 4346 -673
rect -4346 -719 -4238 -685
rect 4238 -719 4346 -685
rect -4346 -731 4346 -719
<< mvnsubdiffcont >>
rect -4238 685 4238 719
rect -4334 -623 -4300 623
rect 4300 -623 4334 623
rect -4238 -719 4238 -685
<< poly >>
rect -4154 581 -4034 597
rect -4154 547 -4138 581
rect -4050 547 -4034 581
rect -4154 500 -4034 547
rect -3976 581 -3856 597
rect -3976 547 -3960 581
rect -3872 547 -3856 581
rect -3976 500 -3856 547
rect -3798 581 -3678 597
rect -3798 547 -3782 581
rect -3694 547 -3678 581
rect -3798 500 -3678 547
rect -3620 581 -3500 597
rect -3620 547 -3604 581
rect -3516 547 -3500 581
rect -3620 500 -3500 547
rect -3442 581 -3322 597
rect -3442 547 -3426 581
rect -3338 547 -3322 581
rect -3442 500 -3322 547
rect -3264 581 -3144 597
rect -3264 547 -3248 581
rect -3160 547 -3144 581
rect -3264 500 -3144 547
rect -3086 581 -2966 597
rect -3086 547 -3070 581
rect -2982 547 -2966 581
rect -3086 500 -2966 547
rect -2908 581 -2788 597
rect -2908 547 -2892 581
rect -2804 547 -2788 581
rect -2908 500 -2788 547
rect -2730 581 -2610 597
rect -2730 547 -2714 581
rect -2626 547 -2610 581
rect -2730 500 -2610 547
rect -2552 581 -2432 597
rect -2552 547 -2536 581
rect -2448 547 -2432 581
rect -2552 500 -2432 547
rect -2374 581 -2254 597
rect -2374 547 -2358 581
rect -2270 547 -2254 581
rect -2374 500 -2254 547
rect -2196 581 -2076 597
rect -2196 547 -2180 581
rect -2092 547 -2076 581
rect -2196 500 -2076 547
rect -2018 581 -1898 597
rect -2018 547 -2002 581
rect -1914 547 -1898 581
rect -2018 500 -1898 547
rect -1840 581 -1720 597
rect -1840 547 -1824 581
rect -1736 547 -1720 581
rect -1840 500 -1720 547
rect -1662 581 -1542 597
rect -1662 547 -1646 581
rect -1558 547 -1542 581
rect -1662 500 -1542 547
rect -1484 581 -1364 597
rect -1484 547 -1468 581
rect -1380 547 -1364 581
rect -1484 500 -1364 547
rect -1306 581 -1186 597
rect -1306 547 -1290 581
rect -1202 547 -1186 581
rect -1306 500 -1186 547
rect -1128 581 -1008 597
rect -1128 547 -1112 581
rect -1024 547 -1008 581
rect -1128 500 -1008 547
rect -950 581 -830 597
rect -950 547 -934 581
rect -846 547 -830 581
rect -950 500 -830 547
rect -772 581 -652 597
rect -772 547 -756 581
rect -668 547 -652 581
rect -772 500 -652 547
rect -594 581 -474 597
rect -594 547 -578 581
rect -490 547 -474 581
rect -594 500 -474 547
rect -416 581 -296 597
rect -416 547 -400 581
rect -312 547 -296 581
rect -416 500 -296 547
rect -238 581 -118 597
rect -238 547 -222 581
rect -134 547 -118 581
rect -238 500 -118 547
rect -60 581 60 597
rect -60 547 -44 581
rect 44 547 60 581
rect -60 500 60 547
rect 118 581 238 597
rect 118 547 134 581
rect 222 547 238 581
rect 118 500 238 547
rect 296 581 416 597
rect 296 547 312 581
rect 400 547 416 581
rect 296 500 416 547
rect 474 581 594 597
rect 474 547 490 581
rect 578 547 594 581
rect 474 500 594 547
rect 652 581 772 597
rect 652 547 668 581
rect 756 547 772 581
rect 652 500 772 547
rect 830 581 950 597
rect 830 547 846 581
rect 934 547 950 581
rect 830 500 950 547
rect 1008 581 1128 597
rect 1008 547 1024 581
rect 1112 547 1128 581
rect 1008 500 1128 547
rect 1186 581 1306 597
rect 1186 547 1202 581
rect 1290 547 1306 581
rect 1186 500 1306 547
rect 1364 581 1484 597
rect 1364 547 1380 581
rect 1468 547 1484 581
rect 1364 500 1484 547
rect 1542 581 1662 597
rect 1542 547 1558 581
rect 1646 547 1662 581
rect 1542 500 1662 547
rect 1720 581 1840 597
rect 1720 547 1736 581
rect 1824 547 1840 581
rect 1720 500 1840 547
rect 1898 581 2018 597
rect 1898 547 1914 581
rect 2002 547 2018 581
rect 1898 500 2018 547
rect 2076 581 2196 597
rect 2076 547 2092 581
rect 2180 547 2196 581
rect 2076 500 2196 547
rect 2254 581 2374 597
rect 2254 547 2270 581
rect 2358 547 2374 581
rect 2254 500 2374 547
rect 2432 581 2552 597
rect 2432 547 2448 581
rect 2536 547 2552 581
rect 2432 500 2552 547
rect 2610 581 2730 597
rect 2610 547 2626 581
rect 2714 547 2730 581
rect 2610 500 2730 547
rect 2788 581 2908 597
rect 2788 547 2804 581
rect 2892 547 2908 581
rect 2788 500 2908 547
rect 2966 581 3086 597
rect 2966 547 2982 581
rect 3070 547 3086 581
rect 2966 500 3086 547
rect 3144 581 3264 597
rect 3144 547 3160 581
rect 3248 547 3264 581
rect 3144 500 3264 547
rect 3322 581 3442 597
rect 3322 547 3338 581
rect 3426 547 3442 581
rect 3322 500 3442 547
rect 3500 581 3620 597
rect 3500 547 3516 581
rect 3604 547 3620 581
rect 3500 500 3620 547
rect 3678 581 3798 597
rect 3678 547 3694 581
rect 3782 547 3798 581
rect 3678 500 3798 547
rect 3856 581 3976 597
rect 3856 547 3872 581
rect 3960 547 3976 581
rect 3856 500 3976 547
rect 4034 581 4154 597
rect 4034 547 4050 581
rect 4138 547 4154 581
rect 4034 500 4154 547
rect -4154 -547 -4034 -500
rect -4154 -581 -4138 -547
rect -4050 -581 -4034 -547
rect -4154 -597 -4034 -581
rect -3976 -547 -3856 -500
rect -3976 -581 -3960 -547
rect -3872 -581 -3856 -547
rect -3976 -597 -3856 -581
rect -3798 -547 -3678 -500
rect -3798 -581 -3782 -547
rect -3694 -581 -3678 -547
rect -3798 -597 -3678 -581
rect -3620 -547 -3500 -500
rect -3620 -581 -3604 -547
rect -3516 -581 -3500 -547
rect -3620 -597 -3500 -581
rect -3442 -547 -3322 -500
rect -3442 -581 -3426 -547
rect -3338 -581 -3322 -547
rect -3442 -597 -3322 -581
rect -3264 -547 -3144 -500
rect -3264 -581 -3248 -547
rect -3160 -581 -3144 -547
rect -3264 -597 -3144 -581
rect -3086 -547 -2966 -500
rect -3086 -581 -3070 -547
rect -2982 -581 -2966 -547
rect -3086 -597 -2966 -581
rect -2908 -547 -2788 -500
rect -2908 -581 -2892 -547
rect -2804 -581 -2788 -547
rect -2908 -597 -2788 -581
rect -2730 -547 -2610 -500
rect -2730 -581 -2714 -547
rect -2626 -581 -2610 -547
rect -2730 -597 -2610 -581
rect -2552 -547 -2432 -500
rect -2552 -581 -2536 -547
rect -2448 -581 -2432 -547
rect -2552 -597 -2432 -581
rect -2374 -547 -2254 -500
rect -2374 -581 -2358 -547
rect -2270 -581 -2254 -547
rect -2374 -597 -2254 -581
rect -2196 -547 -2076 -500
rect -2196 -581 -2180 -547
rect -2092 -581 -2076 -547
rect -2196 -597 -2076 -581
rect -2018 -547 -1898 -500
rect -2018 -581 -2002 -547
rect -1914 -581 -1898 -547
rect -2018 -597 -1898 -581
rect -1840 -547 -1720 -500
rect -1840 -581 -1824 -547
rect -1736 -581 -1720 -547
rect -1840 -597 -1720 -581
rect -1662 -547 -1542 -500
rect -1662 -581 -1646 -547
rect -1558 -581 -1542 -547
rect -1662 -597 -1542 -581
rect -1484 -547 -1364 -500
rect -1484 -581 -1468 -547
rect -1380 -581 -1364 -547
rect -1484 -597 -1364 -581
rect -1306 -547 -1186 -500
rect -1306 -581 -1290 -547
rect -1202 -581 -1186 -547
rect -1306 -597 -1186 -581
rect -1128 -547 -1008 -500
rect -1128 -581 -1112 -547
rect -1024 -581 -1008 -547
rect -1128 -597 -1008 -581
rect -950 -547 -830 -500
rect -950 -581 -934 -547
rect -846 -581 -830 -547
rect -950 -597 -830 -581
rect -772 -547 -652 -500
rect -772 -581 -756 -547
rect -668 -581 -652 -547
rect -772 -597 -652 -581
rect -594 -547 -474 -500
rect -594 -581 -578 -547
rect -490 -581 -474 -547
rect -594 -597 -474 -581
rect -416 -547 -296 -500
rect -416 -581 -400 -547
rect -312 -581 -296 -547
rect -416 -597 -296 -581
rect -238 -547 -118 -500
rect -238 -581 -222 -547
rect -134 -581 -118 -547
rect -238 -597 -118 -581
rect -60 -547 60 -500
rect -60 -581 -44 -547
rect 44 -581 60 -547
rect -60 -597 60 -581
rect 118 -547 238 -500
rect 118 -581 134 -547
rect 222 -581 238 -547
rect 118 -597 238 -581
rect 296 -547 416 -500
rect 296 -581 312 -547
rect 400 -581 416 -547
rect 296 -597 416 -581
rect 474 -547 594 -500
rect 474 -581 490 -547
rect 578 -581 594 -547
rect 474 -597 594 -581
rect 652 -547 772 -500
rect 652 -581 668 -547
rect 756 -581 772 -547
rect 652 -597 772 -581
rect 830 -547 950 -500
rect 830 -581 846 -547
rect 934 -581 950 -547
rect 830 -597 950 -581
rect 1008 -547 1128 -500
rect 1008 -581 1024 -547
rect 1112 -581 1128 -547
rect 1008 -597 1128 -581
rect 1186 -547 1306 -500
rect 1186 -581 1202 -547
rect 1290 -581 1306 -547
rect 1186 -597 1306 -581
rect 1364 -547 1484 -500
rect 1364 -581 1380 -547
rect 1468 -581 1484 -547
rect 1364 -597 1484 -581
rect 1542 -547 1662 -500
rect 1542 -581 1558 -547
rect 1646 -581 1662 -547
rect 1542 -597 1662 -581
rect 1720 -547 1840 -500
rect 1720 -581 1736 -547
rect 1824 -581 1840 -547
rect 1720 -597 1840 -581
rect 1898 -547 2018 -500
rect 1898 -581 1914 -547
rect 2002 -581 2018 -547
rect 1898 -597 2018 -581
rect 2076 -547 2196 -500
rect 2076 -581 2092 -547
rect 2180 -581 2196 -547
rect 2076 -597 2196 -581
rect 2254 -547 2374 -500
rect 2254 -581 2270 -547
rect 2358 -581 2374 -547
rect 2254 -597 2374 -581
rect 2432 -547 2552 -500
rect 2432 -581 2448 -547
rect 2536 -581 2552 -547
rect 2432 -597 2552 -581
rect 2610 -547 2730 -500
rect 2610 -581 2626 -547
rect 2714 -581 2730 -547
rect 2610 -597 2730 -581
rect 2788 -547 2908 -500
rect 2788 -581 2804 -547
rect 2892 -581 2908 -547
rect 2788 -597 2908 -581
rect 2966 -547 3086 -500
rect 2966 -581 2982 -547
rect 3070 -581 3086 -547
rect 2966 -597 3086 -581
rect 3144 -547 3264 -500
rect 3144 -581 3160 -547
rect 3248 -581 3264 -547
rect 3144 -597 3264 -581
rect 3322 -547 3442 -500
rect 3322 -581 3338 -547
rect 3426 -581 3442 -547
rect 3322 -597 3442 -581
rect 3500 -547 3620 -500
rect 3500 -581 3516 -547
rect 3604 -581 3620 -547
rect 3500 -597 3620 -581
rect 3678 -547 3798 -500
rect 3678 -581 3694 -547
rect 3782 -581 3798 -547
rect 3678 -597 3798 -581
rect 3856 -547 3976 -500
rect 3856 -581 3872 -547
rect 3960 -581 3976 -547
rect 3856 -597 3976 -581
rect 4034 -547 4154 -500
rect 4034 -581 4050 -547
rect 4138 -581 4154 -547
rect 4034 -597 4154 -581
<< polycont >>
rect -4138 547 -4050 581
rect -3960 547 -3872 581
rect -3782 547 -3694 581
rect -3604 547 -3516 581
rect -3426 547 -3338 581
rect -3248 547 -3160 581
rect -3070 547 -2982 581
rect -2892 547 -2804 581
rect -2714 547 -2626 581
rect -2536 547 -2448 581
rect -2358 547 -2270 581
rect -2180 547 -2092 581
rect -2002 547 -1914 581
rect -1824 547 -1736 581
rect -1646 547 -1558 581
rect -1468 547 -1380 581
rect -1290 547 -1202 581
rect -1112 547 -1024 581
rect -934 547 -846 581
rect -756 547 -668 581
rect -578 547 -490 581
rect -400 547 -312 581
rect -222 547 -134 581
rect -44 547 44 581
rect 134 547 222 581
rect 312 547 400 581
rect 490 547 578 581
rect 668 547 756 581
rect 846 547 934 581
rect 1024 547 1112 581
rect 1202 547 1290 581
rect 1380 547 1468 581
rect 1558 547 1646 581
rect 1736 547 1824 581
rect 1914 547 2002 581
rect 2092 547 2180 581
rect 2270 547 2358 581
rect 2448 547 2536 581
rect 2626 547 2714 581
rect 2804 547 2892 581
rect 2982 547 3070 581
rect 3160 547 3248 581
rect 3338 547 3426 581
rect 3516 547 3604 581
rect 3694 547 3782 581
rect 3872 547 3960 581
rect 4050 547 4138 581
rect -4138 -581 -4050 -547
rect -3960 -581 -3872 -547
rect -3782 -581 -3694 -547
rect -3604 -581 -3516 -547
rect -3426 -581 -3338 -547
rect -3248 -581 -3160 -547
rect -3070 -581 -2982 -547
rect -2892 -581 -2804 -547
rect -2714 -581 -2626 -547
rect -2536 -581 -2448 -547
rect -2358 -581 -2270 -547
rect -2180 -581 -2092 -547
rect -2002 -581 -1914 -547
rect -1824 -581 -1736 -547
rect -1646 -581 -1558 -547
rect -1468 -581 -1380 -547
rect -1290 -581 -1202 -547
rect -1112 -581 -1024 -547
rect -934 -581 -846 -547
rect -756 -581 -668 -547
rect -578 -581 -490 -547
rect -400 -581 -312 -547
rect -222 -581 -134 -547
rect -44 -581 44 -547
rect 134 -581 222 -547
rect 312 -581 400 -547
rect 490 -581 578 -547
rect 668 -581 756 -547
rect 846 -581 934 -547
rect 1024 -581 1112 -547
rect 1202 -581 1290 -547
rect 1380 -581 1468 -547
rect 1558 -581 1646 -547
rect 1736 -581 1824 -547
rect 1914 -581 2002 -547
rect 2092 -581 2180 -547
rect 2270 -581 2358 -547
rect 2448 -581 2536 -547
rect 2626 -581 2714 -547
rect 2804 -581 2892 -547
rect 2982 -581 3070 -547
rect 3160 -581 3248 -547
rect 3338 -581 3426 -547
rect 3516 -581 3604 -547
rect 3694 -581 3782 -547
rect 3872 -581 3960 -547
rect 4050 -581 4138 -547
<< locali >>
rect -4334 685 -4238 719
rect 4238 685 4334 719
rect -4334 623 -4300 685
rect 4300 623 4334 685
rect -4154 547 -4138 581
rect -4050 547 -4034 581
rect -3976 547 -3960 581
rect -3872 547 -3856 581
rect -3798 547 -3782 581
rect -3694 547 -3678 581
rect -3620 547 -3604 581
rect -3516 547 -3500 581
rect -3442 547 -3426 581
rect -3338 547 -3322 581
rect -3264 547 -3248 581
rect -3160 547 -3144 581
rect -3086 547 -3070 581
rect -2982 547 -2966 581
rect -2908 547 -2892 581
rect -2804 547 -2788 581
rect -2730 547 -2714 581
rect -2626 547 -2610 581
rect -2552 547 -2536 581
rect -2448 547 -2432 581
rect -2374 547 -2358 581
rect -2270 547 -2254 581
rect -2196 547 -2180 581
rect -2092 547 -2076 581
rect -2018 547 -2002 581
rect -1914 547 -1898 581
rect -1840 547 -1824 581
rect -1736 547 -1720 581
rect -1662 547 -1646 581
rect -1558 547 -1542 581
rect -1484 547 -1468 581
rect -1380 547 -1364 581
rect -1306 547 -1290 581
rect -1202 547 -1186 581
rect -1128 547 -1112 581
rect -1024 547 -1008 581
rect -950 547 -934 581
rect -846 547 -830 581
rect -772 547 -756 581
rect -668 547 -652 581
rect -594 547 -578 581
rect -490 547 -474 581
rect -416 547 -400 581
rect -312 547 -296 581
rect -238 547 -222 581
rect -134 547 -118 581
rect -60 547 -44 581
rect 44 547 60 581
rect 118 547 134 581
rect 222 547 238 581
rect 296 547 312 581
rect 400 547 416 581
rect 474 547 490 581
rect 578 547 594 581
rect 652 547 668 581
rect 756 547 772 581
rect 830 547 846 581
rect 934 547 950 581
rect 1008 547 1024 581
rect 1112 547 1128 581
rect 1186 547 1202 581
rect 1290 547 1306 581
rect 1364 547 1380 581
rect 1468 547 1484 581
rect 1542 547 1558 581
rect 1646 547 1662 581
rect 1720 547 1736 581
rect 1824 547 1840 581
rect 1898 547 1914 581
rect 2002 547 2018 581
rect 2076 547 2092 581
rect 2180 547 2196 581
rect 2254 547 2270 581
rect 2358 547 2374 581
rect 2432 547 2448 581
rect 2536 547 2552 581
rect 2610 547 2626 581
rect 2714 547 2730 581
rect 2788 547 2804 581
rect 2892 547 2908 581
rect 2966 547 2982 581
rect 3070 547 3086 581
rect 3144 547 3160 581
rect 3248 547 3264 581
rect 3322 547 3338 581
rect 3426 547 3442 581
rect 3500 547 3516 581
rect 3604 547 3620 581
rect 3678 547 3694 581
rect 3782 547 3798 581
rect 3856 547 3872 581
rect 3960 547 3976 581
rect 4034 547 4050 581
rect 4138 547 4154 581
rect -4200 488 -4166 504
rect -4200 -504 -4166 -488
rect -4022 488 -3988 504
rect -4022 -504 -3988 -488
rect -3844 488 -3810 504
rect -3844 -504 -3810 -488
rect -3666 488 -3632 504
rect -3666 -504 -3632 -488
rect -3488 488 -3454 504
rect -3488 -504 -3454 -488
rect -3310 488 -3276 504
rect -3310 -504 -3276 -488
rect -3132 488 -3098 504
rect -3132 -504 -3098 -488
rect -2954 488 -2920 504
rect -2954 -504 -2920 -488
rect -2776 488 -2742 504
rect -2776 -504 -2742 -488
rect -2598 488 -2564 504
rect -2598 -504 -2564 -488
rect -2420 488 -2386 504
rect -2420 -504 -2386 -488
rect -2242 488 -2208 504
rect -2242 -504 -2208 -488
rect -2064 488 -2030 504
rect -2064 -504 -2030 -488
rect -1886 488 -1852 504
rect -1886 -504 -1852 -488
rect -1708 488 -1674 504
rect -1708 -504 -1674 -488
rect -1530 488 -1496 504
rect -1530 -504 -1496 -488
rect -1352 488 -1318 504
rect -1352 -504 -1318 -488
rect -1174 488 -1140 504
rect -1174 -504 -1140 -488
rect -996 488 -962 504
rect -996 -504 -962 -488
rect -818 488 -784 504
rect -818 -504 -784 -488
rect -640 488 -606 504
rect -640 -504 -606 -488
rect -462 488 -428 504
rect -462 -504 -428 -488
rect -284 488 -250 504
rect -284 -504 -250 -488
rect -106 488 -72 504
rect -106 -504 -72 -488
rect 72 488 106 504
rect 72 -504 106 -488
rect 250 488 284 504
rect 250 -504 284 -488
rect 428 488 462 504
rect 428 -504 462 -488
rect 606 488 640 504
rect 606 -504 640 -488
rect 784 488 818 504
rect 784 -504 818 -488
rect 962 488 996 504
rect 962 -504 996 -488
rect 1140 488 1174 504
rect 1140 -504 1174 -488
rect 1318 488 1352 504
rect 1318 -504 1352 -488
rect 1496 488 1530 504
rect 1496 -504 1530 -488
rect 1674 488 1708 504
rect 1674 -504 1708 -488
rect 1852 488 1886 504
rect 1852 -504 1886 -488
rect 2030 488 2064 504
rect 2030 -504 2064 -488
rect 2208 488 2242 504
rect 2208 -504 2242 -488
rect 2386 488 2420 504
rect 2386 -504 2420 -488
rect 2564 488 2598 504
rect 2564 -504 2598 -488
rect 2742 488 2776 504
rect 2742 -504 2776 -488
rect 2920 488 2954 504
rect 2920 -504 2954 -488
rect 3098 488 3132 504
rect 3098 -504 3132 -488
rect 3276 488 3310 504
rect 3276 -504 3310 -488
rect 3454 488 3488 504
rect 3454 -504 3488 -488
rect 3632 488 3666 504
rect 3632 -504 3666 -488
rect 3810 488 3844 504
rect 3810 -504 3844 -488
rect 3988 488 4022 504
rect 3988 -504 4022 -488
rect 4166 488 4200 504
rect 4166 -504 4200 -488
rect -4154 -581 -4138 -547
rect -4050 -581 -4034 -547
rect -3976 -581 -3960 -547
rect -3872 -581 -3856 -547
rect -3798 -581 -3782 -547
rect -3694 -581 -3678 -547
rect -3620 -581 -3604 -547
rect -3516 -581 -3500 -547
rect -3442 -581 -3426 -547
rect -3338 -581 -3322 -547
rect -3264 -581 -3248 -547
rect -3160 -581 -3144 -547
rect -3086 -581 -3070 -547
rect -2982 -581 -2966 -547
rect -2908 -581 -2892 -547
rect -2804 -581 -2788 -547
rect -2730 -581 -2714 -547
rect -2626 -581 -2610 -547
rect -2552 -581 -2536 -547
rect -2448 -581 -2432 -547
rect -2374 -581 -2358 -547
rect -2270 -581 -2254 -547
rect -2196 -581 -2180 -547
rect -2092 -581 -2076 -547
rect -2018 -581 -2002 -547
rect -1914 -581 -1898 -547
rect -1840 -581 -1824 -547
rect -1736 -581 -1720 -547
rect -1662 -581 -1646 -547
rect -1558 -581 -1542 -547
rect -1484 -581 -1468 -547
rect -1380 -581 -1364 -547
rect -1306 -581 -1290 -547
rect -1202 -581 -1186 -547
rect -1128 -581 -1112 -547
rect -1024 -581 -1008 -547
rect -950 -581 -934 -547
rect -846 -581 -830 -547
rect -772 -581 -756 -547
rect -668 -581 -652 -547
rect -594 -581 -578 -547
rect -490 -581 -474 -547
rect -416 -581 -400 -547
rect -312 -581 -296 -547
rect -238 -581 -222 -547
rect -134 -581 -118 -547
rect -60 -581 -44 -547
rect 44 -581 60 -547
rect 118 -581 134 -547
rect 222 -581 238 -547
rect 296 -581 312 -547
rect 400 -581 416 -547
rect 474 -581 490 -547
rect 578 -581 594 -547
rect 652 -581 668 -547
rect 756 -581 772 -547
rect 830 -581 846 -547
rect 934 -581 950 -547
rect 1008 -581 1024 -547
rect 1112 -581 1128 -547
rect 1186 -581 1202 -547
rect 1290 -581 1306 -547
rect 1364 -581 1380 -547
rect 1468 -581 1484 -547
rect 1542 -581 1558 -547
rect 1646 -581 1662 -547
rect 1720 -581 1736 -547
rect 1824 -581 1840 -547
rect 1898 -581 1914 -547
rect 2002 -581 2018 -547
rect 2076 -581 2092 -547
rect 2180 -581 2196 -547
rect 2254 -581 2270 -547
rect 2358 -581 2374 -547
rect 2432 -581 2448 -547
rect 2536 -581 2552 -547
rect 2610 -581 2626 -547
rect 2714 -581 2730 -547
rect 2788 -581 2804 -547
rect 2892 -581 2908 -547
rect 2966 -581 2982 -547
rect 3070 -581 3086 -547
rect 3144 -581 3160 -547
rect 3248 -581 3264 -547
rect 3322 -581 3338 -547
rect 3426 -581 3442 -547
rect 3500 -581 3516 -547
rect 3604 -581 3620 -547
rect 3678 -581 3694 -547
rect 3782 -581 3798 -547
rect 3856 -581 3872 -547
rect 3960 -581 3976 -547
rect 4034 -581 4050 -547
rect 4138 -581 4154 -547
rect -4334 -685 -4300 -623
rect 4300 -685 4334 -623
rect -4334 -719 -4238 -685
rect 4238 -719 4334 -685
<< viali >>
rect -4138 547 -4050 581
rect -3960 547 -3872 581
rect -3782 547 -3694 581
rect -3604 547 -3516 581
rect -3426 547 -3338 581
rect -3248 547 -3160 581
rect -3070 547 -2982 581
rect -2892 547 -2804 581
rect -2714 547 -2626 581
rect -2536 547 -2448 581
rect -2358 547 -2270 581
rect -2180 547 -2092 581
rect -2002 547 -1914 581
rect -1824 547 -1736 581
rect -1646 547 -1558 581
rect -1468 547 -1380 581
rect -1290 547 -1202 581
rect -1112 547 -1024 581
rect -934 547 -846 581
rect -756 547 -668 581
rect -578 547 -490 581
rect -400 547 -312 581
rect -222 547 -134 581
rect -44 547 44 581
rect 134 547 222 581
rect 312 547 400 581
rect 490 547 578 581
rect 668 547 756 581
rect 846 547 934 581
rect 1024 547 1112 581
rect 1202 547 1290 581
rect 1380 547 1468 581
rect 1558 547 1646 581
rect 1736 547 1824 581
rect 1914 547 2002 581
rect 2092 547 2180 581
rect 2270 547 2358 581
rect 2448 547 2536 581
rect 2626 547 2714 581
rect 2804 547 2892 581
rect 2982 547 3070 581
rect 3160 547 3248 581
rect 3338 547 3426 581
rect 3516 547 3604 581
rect 3694 547 3782 581
rect 3872 547 3960 581
rect 4050 547 4138 581
rect -4200 -488 -4166 488
rect -4022 -488 -3988 488
rect -3844 -488 -3810 488
rect -3666 -488 -3632 488
rect -3488 -488 -3454 488
rect -3310 -488 -3276 488
rect -3132 -488 -3098 488
rect -2954 -488 -2920 488
rect -2776 -488 -2742 488
rect -2598 -488 -2564 488
rect -2420 -488 -2386 488
rect -2242 -488 -2208 488
rect -2064 -488 -2030 488
rect -1886 -488 -1852 488
rect -1708 -488 -1674 488
rect -1530 -488 -1496 488
rect -1352 -488 -1318 488
rect -1174 -488 -1140 488
rect -996 -488 -962 488
rect -818 -488 -784 488
rect -640 -488 -606 488
rect -462 -488 -428 488
rect -284 -488 -250 488
rect -106 -488 -72 488
rect 72 -488 106 488
rect 250 -488 284 488
rect 428 -488 462 488
rect 606 -488 640 488
rect 784 -488 818 488
rect 962 -488 996 488
rect 1140 -488 1174 488
rect 1318 -488 1352 488
rect 1496 -488 1530 488
rect 1674 -488 1708 488
rect 1852 -488 1886 488
rect 2030 -488 2064 488
rect 2208 -488 2242 488
rect 2386 -488 2420 488
rect 2564 -488 2598 488
rect 2742 -488 2776 488
rect 2920 -488 2954 488
rect 3098 -488 3132 488
rect 3276 -488 3310 488
rect 3454 -488 3488 488
rect 3632 -488 3666 488
rect 3810 -488 3844 488
rect 3988 -488 4022 488
rect 4166 -488 4200 488
rect -4138 -581 -4050 -547
rect -3960 -581 -3872 -547
rect -3782 -581 -3694 -547
rect -3604 -581 -3516 -547
rect -3426 -581 -3338 -547
rect -3248 -581 -3160 -547
rect -3070 -581 -2982 -547
rect -2892 -581 -2804 -547
rect -2714 -581 -2626 -547
rect -2536 -581 -2448 -547
rect -2358 -581 -2270 -547
rect -2180 -581 -2092 -547
rect -2002 -581 -1914 -547
rect -1824 -581 -1736 -547
rect -1646 -581 -1558 -547
rect -1468 -581 -1380 -547
rect -1290 -581 -1202 -547
rect -1112 -581 -1024 -547
rect -934 -581 -846 -547
rect -756 -581 -668 -547
rect -578 -581 -490 -547
rect -400 -581 -312 -547
rect -222 -581 -134 -547
rect -44 -581 44 -547
rect 134 -581 222 -547
rect 312 -581 400 -547
rect 490 -581 578 -547
rect 668 -581 756 -547
rect 846 -581 934 -547
rect 1024 -581 1112 -547
rect 1202 -581 1290 -547
rect 1380 -581 1468 -547
rect 1558 -581 1646 -547
rect 1736 -581 1824 -547
rect 1914 -581 2002 -547
rect 2092 -581 2180 -547
rect 2270 -581 2358 -547
rect 2448 -581 2536 -547
rect 2626 -581 2714 -547
rect 2804 -581 2892 -547
rect 2982 -581 3070 -547
rect 3160 -581 3248 -547
rect 3338 -581 3426 -547
rect 3516 -581 3604 -547
rect 3694 -581 3782 -547
rect 3872 -581 3960 -547
rect 4050 -581 4138 -547
<< metal1 >>
rect -4150 581 -4038 587
rect -4150 547 -4138 581
rect -4050 547 -4038 581
rect -4150 541 -4038 547
rect -3972 581 -3860 587
rect -3972 547 -3960 581
rect -3872 547 -3860 581
rect -3972 541 -3860 547
rect -3794 581 -3682 587
rect -3794 547 -3782 581
rect -3694 547 -3682 581
rect -3794 541 -3682 547
rect -3616 581 -3504 587
rect -3616 547 -3604 581
rect -3516 547 -3504 581
rect -3616 541 -3504 547
rect -3438 581 -3326 587
rect -3438 547 -3426 581
rect -3338 547 -3326 581
rect -3438 541 -3326 547
rect -3260 581 -3148 587
rect -3260 547 -3248 581
rect -3160 547 -3148 581
rect -3260 541 -3148 547
rect -3082 581 -2970 587
rect -3082 547 -3070 581
rect -2982 547 -2970 581
rect -3082 541 -2970 547
rect -2904 581 -2792 587
rect -2904 547 -2892 581
rect -2804 547 -2792 581
rect -2904 541 -2792 547
rect -2726 581 -2614 587
rect -2726 547 -2714 581
rect -2626 547 -2614 581
rect -2726 541 -2614 547
rect -2548 581 -2436 587
rect -2548 547 -2536 581
rect -2448 547 -2436 581
rect -2548 541 -2436 547
rect -2370 581 -2258 587
rect -2370 547 -2358 581
rect -2270 547 -2258 581
rect -2370 541 -2258 547
rect -2192 581 -2080 587
rect -2192 547 -2180 581
rect -2092 547 -2080 581
rect -2192 541 -2080 547
rect -2014 581 -1902 587
rect -2014 547 -2002 581
rect -1914 547 -1902 581
rect -2014 541 -1902 547
rect -1836 581 -1724 587
rect -1836 547 -1824 581
rect -1736 547 -1724 581
rect -1836 541 -1724 547
rect -1658 581 -1546 587
rect -1658 547 -1646 581
rect -1558 547 -1546 581
rect -1658 541 -1546 547
rect -1480 581 -1368 587
rect -1480 547 -1468 581
rect -1380 547 -1368 581
rect -1480 541 -1368 547
rect -1302 581 -1190 587
rect -1302 547 -1290 581
rect -1202 547 -1190 581
rect -1302 541 -1190 547
rect -1124 581 -1012 587
rect -1124 547 -1112 581
rect -1024 547 -1012 581
rect -1124 541 -1012 547
rect -946 581 -834 587
rect -946 547 -934 581
rect -846 547 -834 581
rect -946 541 -834 547
rect -768 581 -656 587
rect -768 547 -756 581
rect -668 547 -656 581
rect -768 541 -656 547
rect -590 581 -478 587
rect -590 547 -578 581
rect -490 547 -478 581
rect -590 541 -478 547
rect -412 581 -300 587
rect -412 547 -400 581
rect -312 547 -300 581
rect -412 541 -300 547
rect -234 581 -122 587
rect -234 547 -222 581
rect -134 547 -122 581
rect -234 541 -122 547
rect -56 581 56 587
rect -56 547 -44 581
rect 44 547 56 581
rect -56 541 56 547
rect 122 581 234 587
rect 122 547 134 581
rect 222 547 234 581
rect 122 541 234 547
rect 300 581 412 587
rect 300 547 312 581
rect 400 547 412 581
rect 300 541 412 547
rect 478 581 590 587
rect 478 547 490 581
rect 578 547 590 581
rect 478 541 590 547
rect 656 581 768 587
rect 656 547 668 581
rect 756 547 768 581
rect 656 541 768 547
rect 834 581 946 587
rect 834 547 846 581
rect 934 547 946 581
rect 834 541 946 547
rect 1012 581 1124 587
rect 1012 547 1024 581
rect 1112 547 1124 581
rect 1012 541 1124 547
rect 1190 581 1302 587
rect 1190 547 1202 581
rect 1290 547 1302 581
rect 1190 541 1302 547
rect 1368 581 1480 587
rect 1368 547 1380 581
rect 1468 547 1480 581
rect 1368 541 1480 547
rect 1546 581 1658 587
rect 1546 547 1558 581
rect 1646 547 1658 581
rect 1546 541 1658 547
rect 1724 581 1836 587
rect 1724 547 1736 581
rect 1824 547 1836 581
rect 1724 541 1836 547
rect 1902 581 2014 587
rect 1902 547 1914 581
rect 2002 547 2014 581
rect 1902 541 2014 547
rect 2080 581 2192 587
rect 2080 547 2092 581
rect 2180 547 2192 581
rect 2080 541 2192 547
rect 2258 581 2370 587
rect 2258 547 2270 581
rect 2358 547 2370 581
rect 2258 541 2370 547
rect 2436 581 2548 587
rect 2436 547 2448 581
rect 2536 547 2548 581
rect 2436 541 2548 547
rect 2614 581 2726 587
rect 2614 547 2626 581
rect 2714 547 2726 581
rect 2614 541 2726 547
rect 2792 581 2904 587
rect 2792 547 2804 581
rect 2892 547 2904 581
rect 2792 541 2904 547
rect 2970 581 3082 587
rect 2970 547 2982 581
rect 3070 547 3082 581
rect 2970 541 3082 547
rect 3148 581 3260 587
rect 3148 547 3160 581
rect 3248 547 3260 581
rect 3148 541 3260 547
rect 3326 581 3438 587
rect 3326 547 3338 581
rect 3426 547 3438 581
rect 3326 541 3438 547
rect 3504 581 3616 587
rect 3504 547 3516 581
rect 3604 547 3616 581
rect 3504 541 3616 547
rect 3682 581 3794 587
rect 3682 547 3694 581
rect 3782 547 3794 581
rect 3682 541 3794 547
rect 3860 581 3972 587
rect 3860 547 3872 581
rect 3960 547 3972 581
rect 3860 541 3972 547
rect 4038 581 4150 587
rect 4038 547 4050 581
rect 4138 547 4150 581
rect 4038 541 4150 547
rect -4206 488 -4160 500
rect -4206 -488 -4200 488
rect -4166 -488 -4160 488
rect -4206 -500 -4160 -488
rect -4028 488 -3982 500
rect -4028 -488 -4022 488
rect -3988 -488 -3982 488
rect -4028 -500 -3982 -488
rect -3850 488 -3804 500
rect -3850 -488 -3844 488
rect -3810 -488 -3804 488
rect -3850 -500 -3804 -488
rect -3672 488 -3626 500
rect -3672 -488 -3666 488
rect -3632 -488 -3626 488
rect -3672 -500 -3626 -488
rect -3494 488 -3448 500
rect -3494 -488 -3488 488
rect -3454 -488 -3448 488
rect -3494 -500 -3448 -488
rect -3316 488 -3270 500
rect -3316 -488 -3310 488
rect -3276 -488 -3270 488
rect -3316 -500 -3270 -488
rect -3138 488 -3092 500
rect -3138 -488 -3132 488
rect -3098 -488 -3092 488
rect -3138 -500 -3092 -488
rect -2960 488 -2914 500
rect -2960 -488 -2954 488
rect -2920 -488 -2914 488
rect -2960 -500 -2914 -488
rect -2782 488 -2736 500
rect -2782 -488 -2776 488
rect -2742 -488 -2736 488
rect -2782 -500 -2736 -488
rect -2604 488 -2558 500
rect -2604 -488 -2598 488
rect -2564 -488 -2558 488
rect -2604 -500 -2558 -488
rect -2426 488 -2380 500
rect -2426 -488 -2420 488
rect -2386 -488 -2380 488
rect -2426 -500 -2380 -488
rect -2248 488 -2202 500
rect -2248 -488 -2242 488
rect -2208 -488 -2202 488
rect -2248 -500 -2202 -488
rect -2070 488 -2024 500
rect -2070 -488 -2064 488
rect -2030 -488 -2024 488
rect -2070 -500 -2024 -488
rect -1892 488 -1846 500
rect -1892 -488 -1886 488
rect -1852 -488 -1846 488
rect -1892 -500 -1846 -488
rect -1714 488 -1668 500
rect -1714 -488 -1708 488
rect -1674 -488 -1668 488
rect -1714 -500 -1668 -488
rect -1536 488 -1490 500
rect -1536 -488 -1530 488
rect -1496 -488 -1490 488
rect -1536 -500 -1490 -488
rect -1358 488 -1312 500
rect -1358 -488 -1352 488
rect -1318 -488 -1312 488
rect -1358 -500 -1312 -488
rect -1180 488 -1134 500
rect -1180 -488 -1174 488
rect -1140 -488 -1134 488
rect -1180 -500 -1134 -488
rect -1002 488 -956 500
rect -1002 -488 -996 488
rect -962 -488 -956 488
rect -1002 -500 -956 -488
rect -824 488 -778 500
rect -824 -488 -818 488
rect -784 -488 -778 488
rect -824 -500 -778 -488
rect -646 488 -600 500
rect -646 -488 -640 488
rect -606 -488 -600 488
rect -646 -500 -600 -488
rect -468 488 -422 500
rect -468 -488 -462 488
rect -428 -488 -422 488
rect -468 -500 -422 -488
rect -290 488 -244 500
rect -290 -488 -284 488
rect -250 -488 -244 488
rect -290 -500 -244 -488
rect -112 488 -66 500
rect -112 -488 -106 488
rect -72 -488 -66 488
rect -112 -500 -66 -488
rect 66 488 112 500
rect 66 -488 72 488
rect 106 -488 112 488
rect 66 -500 112 -488
rect 244 488 290 500
rect 244 -488 250 488
rect 284 -488 290 488
rect 244 -500 290 -488
rect 422 488 468 500
rect 422 -488 428 488
rect 462 -488 468 488
rect 422 -500 468 -488
rect 600 488 646 500
rect 600 -488 606 488
rect 640 -488 646 488
rect 600 -500 646 -488
rect 778 488 824 500
rect 778 -488 784 488
rect 818 -488 824 488
rect 778 -500 824 -488
rect 956 488 1002 500
rect 956 -488 962 488
rect 996 -488 1002 488
rect 956 -500 1002 -488
rect 1134 488 1180 500
rect 1134 -488 1140 488
rect 1174 -488 1180 488
rect 1134 -500 1180 -488
rect 1312 488 1358 500
rect 1312 -488 1318 488
rect 1352 -488 1358 488
rect 1312 -500 1358 -488
rect 1490 488 1536 500
rect 1490 -488 1496 488
rect 1530 -488 1536 488
rect 1490 -500 1536 -488
rect 1668 488 1714 500
rect 1668 -488 1674 488
rect 1708 -488 1714 488
rect 1668 -500 1714 -488
rect 1846 488 1892 500
rect 1846 -488 1852 488
rect 1886 -488 1892 488
rect 1846 -500 1892 -488
rect 2024 488 2070 500
rect 2024 -488 2030 488
rect 2064 -488 2070 488
rect 2024 -500 2070 -488
rect 2202 488 2248 500
rect 2202 -488 2208 488
rect 2242 -488 2248 488
rect 2202 -500 2248 -488
rect 2380 488 2426 500
rect 2380 -488 2386 488
rect 2420 -488 2426 488
rect 2380 -500 2426 -488
rect 2558 488 2604 500
rect 2558 -488 2564 488
rect 2598 -488 2604 488
rect 2558 -500 2604 -488
rect 2736 488 2782 500
rect 2736 -488 2742 488
rect 2776 -488 2782 488
rect 2736 -500 2782 -488
rect 2914 488 2960 500
rect 2914 -488 2920 488
rect 2954 -488 2960 488
rect 2914 -500 2960 -488
rect 3092 488 3138 500
rect 3092 -488 3098 488
rect 3132 -488 3138 488
rect 3092 -500 3138 -488
rect 3270 488 3316 500
rect 3270 -488 3276 488
rect 3310 -488 3316 488
rect 3270 -500 3316 -488
rect 3448 488 3494 500
rect 3448 -488 3454 488
rect 3488 -488 3494 488
rect 3448 -500 3494 -488
rect 3626 488 3672 500
rect 3626 -488 3632 488
rect 3666 -488 3672 488
rect 3626 -500 3672 -488
rect 3804 488 3850 500
rect 3804 -488 3810 488
rect 3844 -488 3850 488
rect 3804 -500 3850 -488
rect 3982 488 4028 500
rect 3982 -488 3988 488
rect 4022 -488 4028 488
rect 3982 -500 4028 -488
rect 4160 488 4206 500
rect 4160 -488 4166 488
rect 4200 -488 4206 488
rect 4160 -500 4206 -488
rect -4150 -547 -4038 -541
rect -4150 -581 -4138 -547
rect -4050 -581 -4038 -547
rect -4150 -587 -4038 -581
rect -3972 -547 -3860 -541
rect -3972 -581 -3960 -547
rect -3872 -581 -3860 -547
rect -3972 -587 -3860 -581
rect -3794 -547 -3682 -541
rect -3794 -581 -3782 -547
rect -3694 -581 -3682 -547
rect -3794 -587 -3682 -581
rect -3616 -547 -3504 -541
rect -3616 -581 -3604 -547
rect -3516 -581 -3504 -547
rect -3616 -587 -3504 -581
rect -3438 -547 -3326 -541
rect -3438 -581 -3426 -547
rect -3338 -581 -3326 -547
rect -3438 -587 -3326 -581
rect -3260 -547 -3148 -541
rect -3260 -581 -3248 -547
rect -3160 -581 -3148 -547
rect -3260 -587 -3148 -581
rect -3082 -547 -2970 -541
rect -3082 -581 -3070 -547
rect -2982 -581 -2970 -547
rect -3082 -587 -2970 -581
rect -2904 -547 -2792 -541
rect -2904 -581 -2892 -547
rect -2804 -581 -2792 -547
rect -2904 -587 -2792 -581
rect -2726 -547 -2614 -541
rect -2726 -581 -2714 -547
rect -2626 -581 -2614 -547
rect -2726 -587 -2614 -581
rect -2548 -547 -2436 -541
rect -2548 -581 -2536 -547
rect -2448 -581 -2436 -547
rect -2548 -587 -2436 -581
rect -2370 -547 -2258 -541
rect -2370 -581 -2358 -547
rect -2270 -581 -2258 -547
rect -2370 -587 -2258 -581
rect -2192 -547 -2080 -541
rect -2192 -581 -2180 -547
rect -2092 -581 -2080 -547
rect -2192 -587 -2080 -581
rect -2014 -547 -1902 -541
rect -2014 -581 -2002 -547
rect -1914 -581 -1902 -547
rect -2014 -587 -1902 -581
rect -1836 -547 -1724 -541
rect -1836 -581 -1824 -547
rect -1736 -581 -1724 -547
rect -1836 -587 -1724 -581
rect -1658 -547 -1546 -541
rect -1658 -581 -1646 -547
rect -1558 -581 -1546 -547
rect -1658 -587 -1546 -581
rect -1480 -547 -1368 -541
rect -1480 -581 -1468 -547
rect -1380 -581 -1368 -547
rect -1480 -587 -1368 -581
rect -1302 -547 -1190 -541
rect -1302 -581 -1290 -547
rect -1202 -581 -1190 -547
rect -1302 -587 -1190 -581
rect -1124 -547 -1012 -541
rect -1124 -581 -1112 -547
rect -1024 -581 -1012 -547
rect -1124 -587 -1012 -581
rect -946 -547 -834 -541
rect -946 -581 -934 -547
rect -846 -581 -834 -547
rect -946 -587 -834 -581
rect -768 -547 -656 -541
rect -768 -581 -756 -547
rect -668 -581 -656 -547
rect -768 -587 -656 -581
rect -590 -547 -478 -541
rect -590 -581 -578 -547
rect -490 -581 -478 -547
rect -590 -587 -478 -581
rect -412 -547 -300 -541
rect -412 -581 -400 -547
rect -312 -581 -300 -547
rect -412 -587 -300 -581
rect -234 -547 -122 -541
rect -234 -581 -222 -547
rect -134 -581 -122 -547
rect -234 -587 -122 -581
rect -56 -547 56 -541
rect -56 -581 -44 -547
rect 44 -581 56 -547
rect -56 -587 56 -581
rect 122 -547 234 -541
rect 122 -581 134 -547
rect 222 -581 234 -547
rect 122 -587 234 -581
rect 300 -547 412 -541
rect 300 -581 312 -547
rect 400 -581 412 -547
rect 300 -587 412 -581
rect 478 -547 590 -541
rect 478 -581 490 -547
rect 578 -581 590 -547
rect 478 -587 590 -581
rect 656 -547 768 -541
rect 656 -581 668 -547
rect 756 -581 768 -547
rect 656 -587 768 -581
rect 834 -547 946 -541
rect 834 -581 846 -547
rect 934 -581 946 -547
rect 834 -587 946 -581
rect 1012 -547 1124 -541
rect 1012 -581 1024 -547
rect 1112 -581 1124 -547
rect 1012 -587 1124 -581
rect 1190 -547 1302 -541
rect 1190 -581 1202 -547
rect 1290 -581 1302 -547
rect 1190 -587 1302 -581
rect 1368 -547 1480 -541
rect 1368 -581 1380 -547
rect 1468 -581 1480 -547
rect 1368 -587 1480 -581
rect 1546 -547 1658 -541
rect 1546 -581 1558 -547
rect 1646 -581 1658 -547
rect 1546 -587 1658 -581
rect 1724 -547 1836 -541
rect 1724 -581 1736 -547
rect 1824 -581 1836 -547
rect 1724 -587 1836 -581
rect 1902 -547 2014 -541
rect 1902 -581 1914 -547
rect 2002 -581 2014 -547
rect 1902 -587 2014 -581
rect 2080 -547 2192 -541
rect 2080 -581 2092 -547
rect 2180 -581 2192 -547
rect 2080 -587 2192 -581
rect 2258 -547 2370 -541
rect 2258 -581 2270 -547
rect 2358 -581 2370 -547
rect 2258 -587 2370 -581
rect 2436 -547 2548 -541
rect 2436 -581 2448 -547
rect 2536 -581 2548 -547
rect 2436 -587 2548 -581
rect 2614 -547 2726 -541
rect 2614 -581 2626 -547
rect 2714 -581 2726 -547
rect 2614 -587 2726 -581
rect 2792 -547 2904 -541
rect 2792 -581 2804 -547
rect 2892 -581 2904 -547
rect 2792 -587 2904 -581
rect 2970 -547 3082 -541
rect 2970 -581 2982 -547
rect 3070 -581 3082 -547
rect 2970 -587 3082 -581
rect 3148 -547 3260 -541
rect 3148 -581 3160 -547
rect 3248 -581 3260 -547
rect 3148 -587 3260 -581
rect 3326 -547 3438 -541
rect 3326 -581 3338 -547
rect 3426 -581 3438 -547
rect 3326 -587 3438 -581
rect 3504 -547 3616 -541
rect 3504 -581 3516 -547
rect 3604 -581 3616 -547
rect 3504 -587 3616 -581
rect 3682 -547 3794 -541
rect 3682 -581 3694 -547
rect 3782 -581 3794 -547
rect 3682 -587 3794 -581
rect 3860 -547 3972 -541
rect 3860 -581 3872 -547
rect 3960 -581 3972 -547
rect 3860 -587 3972 -581
rect 4038 -547 4150 -541
rect 4038 -581 4050 -547
rect 4138 -581 4150 -547
rect 4038 -587 4150 -581
<< properties >>
string FIXED_BBOX -4317 -702 4317 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.6 m 1 nf 47 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
