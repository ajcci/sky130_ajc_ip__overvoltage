** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/comparator_wip.sch
**.subckt comparator_wip ena avdd avss ibias vinn vinp out
*.ipin ena
*.ipin avdd
*.ipin avss
*.ipin ibias
*.ipin vinn
*.ipin vinp
*.opin out
XMi0 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8e-06 W=4.2e-07 m=16 
XMi1 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8e-06 W=4.2e-07 m=16 
XMb vn vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8e-06 W=1e-06 m=2 
XMta vt vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8e-06 W=1e-06 m=2 
XMld1 vpp vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8e-06 W=4.2e-07 m=8 
XMh1 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8e-06 W=4.2e-07 m=10 
XMh0 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8e-06 W=4.2e-07 m=10 
XMld0 vnn vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8e-06 W=4.2e-07 m=8 
XMnn1 n0 vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8e-06 W=1e-06 m=2 
XMnn0 vm vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8e-06 W=1e-06 m=2 
XMpp1 n0 vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8e-06 W=1e-06 m=2 
XMpp0 vm vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8e-06 W=1e-06 m=2 
**.ends
.end
