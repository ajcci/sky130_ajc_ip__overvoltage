magic
tech sky130A
timestamp 1712158818
<< pwell >>
rect -2191 -379 2191 379
<< mvnmos >>
rect -2077 -250 -2017 250
rect -1988 -250 -1928 250
rect -1899 -250 -1839 250
rect -1810 -250 -1750 250
rect -1721 -250 -1661 250
rect -1632 -250 -1572 250
rect -1543 -250 -1483 250
rect -1454 -250 -1394 250
rect -1365 -250 -1305 250
rect -1276 -250 -1216 250
rect -1187 -250 -1127 250
rect -1098 -250 -1038 250
rect -1009 -250 -949 250
rect -920 -250 -860 250
rect -831 -250 -771 250
rect -742 -250 -682 250
rect -653 -250 -593 250
rect -564 -250 -504 250
rect -475 -250 -415 250
rect -386 -250 -326 250
rect -297 -250 -237 250
rect -208 -250 -148 250
rect -119 -250 -59 250
rect -30 -250 30 250
rect 59 -250 119 250
rect 148 -250 208 250
rect 237 -250 297 250
rect 326 -250 386 250
rect 415 -250 475 250
rect 504 -250 564 250
rect 593 -250 653 250
rect 682 -250 742 250
rect 771 -250 831 250
rect 860 -250 920 250
rect 949 -250 1009 250
rect 1038 -250 1098 250
rect 1127 -250 1187 250
rect 1216 -250 1276 250
rect 1305 -250 1365 250
rect 1394 -250 1454 250
rect 1483 -250 1543 250
rect 1572 -250 1632 250
rect 1661 -250 1721 250
rect 1750 -250 1810 250
rect 1839 -250 1899 250
rect 1928 -250 1988 250
rect 2017 -250 2077 250
<< mvndiff >>
rect -2106 244 -2077 250
rect -2106 -244 -2100 244
rect -2083 -244 -2077 244
rect -2106 -250 -2077 -244
rect -2017 244 -1988 250
rect -2017 -244 -2011 244
rect -1994 -244 -1988 244
rect -2017 -250 -1988 -244
rect -1928 244 -1899 250
rect -1928 -244 -1922 244
rect -1905 -244 -1899 244
rect -1928 -250 -1899 -244
rect -1839 244 -1810 250
rect -1839 -244 -1833 244
rect -1816 -244 -1810 244
rect -1839 -250 -1810 -244
rect -1750 244 -1721 250
rect -1750 -244 -1744 244
rect -1727 -244 -1721 244
rect -1750 -250 -1721 -244
rect -1661 244 -1632 250
rect -1661 -244 -1655 244
rect -1638 -244 -1632 244
rect -1661 -250 -1632 -244
rect -1572 244 -1543 250
rect -1572 -244 -1566 244
rect -1549 -244 -1543 244
rect -1572 -250 -1543 -244
rect -1483 244 -1454 250
rect -1483 -244 -1477 244
rect -1460 -244 -1454 244
rect -1483 -250 -1454 -244
rect -1394 244 -1365 250
rect -1394 -244 -1388 244
rect -1371 -244 -1365 244
rect -1394 -250 -1365 -244
rect -1305 244 -1276 250
rect -1305 -244 -1299 244
rect -1282 -244 -1276 244
rect -1305 -250 -1276 -244
rect -1216 244 -1187 250
rect -1216 -244 -1210 244
rect -1193 -244 -1187 244
rect -1216 -250 -1187 -244
rect -1127 244 -1098 250
rect -1127 -244 -1121 244
rect -1104 -244 -1098 244
rect -1127 -250 -1098 -244
rect -1038 244 -1009 250
rect -1038 -244 -1032 244
rect -1015 -244 -1009 244
rect -1038 -250 -1009 -244
rect -949 244 -920 250
rect -949 -244 -943 244
rect -926 -244 -920 244
rect -949 -250 -920 -244
rect -860 244 -831 250
rect -860 -244 -854 244
rect -837 -244 -831 244
rect -860 -250 -831 -244
rect -771 244 -742 250
rect -771 -244 -765 244
rect -748 -244 -742 244
rect -771 -250 -742 -244
rect -682 244 -653 250
rect -682 -244 -676 244
rect -659 -244 -653 244
rect -682 -250 -653 -244
rect -593 244 -564 250
rect -593 -244 -587 244
rect -570 -244 -564 244
rect -593 -250 -564 -244
rect -504 244 -475 250
rect -504 -244 -498 244
rect -481 -244 -475 244
rect -504 -250 -475 -244
rect -415 244 -386 250
rect -415 -244 -409 244
rect -392 -244 -386 244
rect -415 -250 -386 -244
rect -326 244 -297 250
rect -326 -244 -320 244
rect -303 -244 -297 244
rect -326 -250 -297 -244
rect -237 244 -208 250
rect -237 -244 -231 244
rect -214 -244 -208 244
rect -237 -250 -208 -244
rect -148 244 -119 250
rect -148 -244 -142 244
rect -125 -244 -119 244
rect -148 -250 -119 -244
rect -59 244 -30 250
rect -59 -244 -53 244
rect -36 -244 -30 244
rect -59 -250 -30 -244
rect 30 244 59 250
rect 30 -244 36 244
rect 53 -244 59 244
rect 30 -250 59 -244
rect 119 244 148 250
rect 119 -244 125 244
rect 142 -244 148 244
rect 119 -250 148 -244
rect 208 244 237 250
rect 208 -244 214 244
rect 231 -244 237 244
rect 208 -250 237 -244
rect 297 244 326 250
rect 297 -244 303 244
rect 320 -244 326 244
rect 297 -250 326 -244
rect 386 244 415 250
rect 386 -244 392 244
rect 409 -244 415 244
rect 386 -250 415 -244
rect 475 244 504 250
rect 475 -244 481 244
rect 498 -244 504 244
rect 475 -250 504 -244
rect 564 244 593 250
rect 564 -244 570 244
rect 587 -244 593 244
rect 564 -250 593 -244
rect 653 244 682 250
rect 653 -244 659 244
rect 676 -244 682 244
rect 653 -250 682 -244
rect 742 244 771 250
rect 742 -244 748 244
rect 765 -244 771 244
rect 742 -250 771 -244
rect 831 244 860 250
rect 831 -244 837 244
rect 854 -244 860 244
rect 831 -250 860 -244
rect 920 244 949 250
rect 920 -244 926 244
rect 943 -244 949 244
rect 920 -250 949 -244
rect 1009 244 1038 250
rect 1009 -244 1015 244
rect 1032 -244 1038 244
rect 1009 -250 1038 -244
rect 1098 244 1127 250
rect 1098 -244 1104 244
rect 1121 -244 1127 244
rect 1098 -250 1127 -244
rect 1187 244 1216 250
rect 1187 -244 1193 244
rect 1210 -244 1216 244
rect 1187 -250 1216 -244
rect 1276 244 1305 250
rect 1276 -244 1282 244
rect 1299 -244 1305 244
rect 1276 -250 1305 -244
rect 1365 244 1394 250
rect 1365 -244 1371 244
rect 1388 -244 1394 244
rect 1365 -250 1394 -244
rect 1454 244 1483 250
rect 1454 -244 1460 244
rect 1477 -244 1483 244
rect 1454 -250 1483 -244
rect 1543 244 1572 250
rect 1543 -244 1549 244
rect 1566 -244 1572 244
rect 1543 -250 1572 -244
rect 1632 244 1661 250
rect 1632 -244 1638 244
rect 1655 -244 1661 244
rect 1632 -250 1661 -244
rect 1721 244 1750 250
rect 1721 -244 1727 244
rect 1744 -244 1750 244
rect 1721 -250 1750 -244
rect 1810 244 1839 250
rect 1810 -244 1816 244
rect 1833 -244 1839 244
rect 1810 -250 1839 -244
rect 1899 244 1928 250
rect 1899 -244 1905 244
rect 1922 -244 1928 244
rect 1899 -250 1928 -244
rect 1988 244 2017 250
rect 1988 -244 1994 244
rect 2011 -244 2017 244
rect 1988 -250 2017 -244
rect 2077 244 2106 250
rect 2077 -244 2083 244
rect 2100 -244 2106 244
rect 2077 -250 2106 -244
<< mvndiffc >>
rect -2100 -244 -2083 244
rect -2011 -244 -1994 244
rect -1922 -244 -1905 244
rect -1833 -244 -1816 244
rect -1744 -244 -1727 244
rect -1655 -244 -1638 244
rect -1566 -244 -1549 244
rect -1477 -244 -1460 244
rect -1388 -244 -1371 244
rect -1299 -244 -1282 244
rect -1210 -244 -1193 244
rect -1121 -244 -1104 244
rect -1032 -244 -1015 244
rect -943 -244 -926 244
rect -854 -244 -837 244
rect -765 -244 -748 244
rect -676 -244 -659 244
rect -587 -244 -570 244
rect -498 -244 -481 244
rect -409 -244 -392 244
rect -320 -244 -303 244
rect -231 -244 -214 244
rect -142 -244 -125 244
rect -53 -244 -36 244
rect 36 -244 53 244
rect 125 -244 142 244
rect 214 -244 231 244
rect 303 -244 320 244
rect 392 -244 409 244
rect 481 -244 498 244
rect 570 -244 587 244
rect 659 -244 676 244
rect 748 -244 765 244
rect 837 -244 854 244
rect 926 -244 943 244
rect 1015 -244 1032 244
rect 1104 -244 1121 244
rect 1193 -244 1210 244
rect 1282 -244 1299 244
rect 1371 -244 1388 244
rect 1460 -244 1477 244
rect 1549 -244 1566 244
rect 1638 -244 1655 244
rect 1727 -244 1744 244
rect 1816 -244 1833 244
rect 1905 -244 1922 244
rect 1994 -244 2011 244
rect 2083 -244 2100 244
<< mvpsubdiff >>
rect -2173 355 2173 361
rect -2173 338 -2119 355
rect 2119 338 2173 355
rect -2173 332 2173 338
rect -2173 307 -2144 332
rect -2173 -307 -2167 307
rect -2150 -307 -2144 307
rect 2144 307 2173 332
rect -2173 -332 -2144 -307
rect 2144 -307 2150 307
rect 2167 -307 2173 307
rect 2144 -332 2173 -307
rect -2173 -338 2173 -332
rect -2173 -355 -2119 -338
rect 2119 -355 2173 -338
rect -2173 -361 2173 -355
<< mvpsubdiffcont >>
rect -2119 338 2119 355
rect -2167 -307 -2150 307
rect 2150 -307 2167 307
rect -2119 -355 2119 -338
<< poly >>
rect -2077 286 -2017 294
rect -2077 269 -2069 286
rect -2025 269 -2017 286
rect -2077 250 -2017 269
rect -1988 286 -1928 294
rect -1988 269 -1980 286
rect -1936 269 -1928 286
rect -1988 250 -1928 269
rect -1899 286 -1839 294
rect -1899 269 -1891 286
rect -1847 269 -1839 286
rect -1899 250 -1839 269
rect -1810 286 -1750 294
rect -1810 269 -1802 286
rect -1758 269 -1750 286
rect -1810 250 -1750 269
rect -1721 286 -1661 294
rect -1721 269 -1713 286
rect -1669 269 -1661 286
rect -1721 250 -1661 269
rect -1632 286 -1572 294
rect -1632 269 -1624 286
rect -1580 269 -1572 286
rect -1632 250 -1572 269
rect -1543 286 -1483 294
rect -1543 269 -1535 286
rect -1491 269 -1483 286
rect -1543 250 -1483 269
rect -1454 286 -1394 294
rect -1454 269 -1446 286
rect -1402 269 -1394 286
rect -1454 250 -1394 269
rect -1365 286 -1305 294
rect -1365 269 -1357 286
rect -1313 269 -1305 286
rect -1365 250 -1305 269
rect -1276 286 -1216 294
rect -1276 269 -1268 286
rect -1224 269 -1216 286
rect -1276 250 -1216 269
rect -1187 286 -1127 294
rect -1187 269 -1179 286
rect -1135 269 -1127 286
rect -1187 250 -1127 269
rect -1098 286 -1038 294
rect -1098 269 -1090 286
rect -1046 269 -1038 286
rect -1098 250 -1038 269
rect -1009 286 -949 294
rect -1009 269 -1001 286
rect -957 269 -949 286
rect -1009 250 -949 269
rect -920 286 -860 294
rect -920 269 -912 286
rect -868 269 -860 286
rect -920 250 -860 269
rect -831 286 -771 294
rect -831 269 -823 286
rect -779 269 -771 286
rect -831 250 -771 269
rect -742 286 -682 294
rect -742 269 -734 286
rect -690 269 -682 286
rect -742 250 -682 269
rect -653 286 -593 294
rect -653 269 -645 286
rect -601 269 -593 286
rect -653 250 -593 269
rect -564 286 -504 294
rect -564 269 -556 286
rect -512 269 -504 286
rect -564 250 -504 269
rect -475 286 -415 294
rect -475 269 -467 286
rect -423 269 -415 286
rect -475 250 -415 269
rect -386 286 -326 294
rect -386 269 -378 286
rect -334 269 -326 286
rect -386 250 -326 269
rect -297 286 -237 294
rect -297 269 -289 286
rect -245 269 -237 286
rect -297 250 -237 269
rect -208 286 -148 294
rect -208 269 -200 286
rect -156 269 -148 286
rect -208 250 -148 269
rect -119 286 -59 294
rect -119 269 -111 286
rect -67 269 -59 286
rect -119 250 -59 269
rect -30 286 30 294
rect -30 269 -22 286
rect 22 269 30 286
rect -30 250 30 269
rect 59 286 119 294
rect 59 269 67 286
rect 111 269 119 286
rect 59 250 119 269
rect 148 286 208 294
rect 148 269 156 286
rect 200 269 208 286
rect 148 250 208 269
rect 237 286 297 294
rect 237 269 245 286
rect 289 269 297 286
rect 237 250 297 269
rect 326 286 386 294
rect 326 269 334 286
rect 378 269 386 286
rect 326 250 386 269
rect 415 286 475 294
rect 415 269 423 286
rect 467 269 475 286
rect 415 250 475 269
rect 504 286 564 294
rect 504 269 512 286
rect 556 269 564 286
rect 504 250 564 269
rect 593 286 653 294
rect 593 269 601 286
rect 645 269 653 286
rect 593 250 653 269
rect 682 286 742 294
rect 682 269 690 286
rect 734 269 742 286
rect 682 250 742 269
rect 771 286 831 294
rect 771 269 779 286
rect 823 269 831 286
rect 771 250 831 269
rect 860 286 920 294
rect 860 269 868 286
rect 912 269 920 286
rect 860 250 920 269
rect 949 286 1009 294
rect 949 269 957 286
rect 1001 269 1009 286
rect 949 250 1009 269
rect 1038 286 1098 294
rect 1038 269 1046 286
rect 1090 269 1098 286
rect 1038 250 1098 269
rect 1127 286 1187 294
rect 1127 269 1135 286
rect 1179 269 1187 286
rect 1127 250 1187 269
rect 1216 286 1276 294
rect 1216 269 1224 286
rect 1268 269 1276 286
rect 1216 250 1276 269
rect 1305 286 1365 294
rect 1305 269 1313 286
rect 1357 269 1365 286
rect 1305 250 1365 269
rect 1394 286 1454 294
rect 1394 269 1402 286
rect 1446 269 1454 286
rect 1394 250 1454 269
rect 1483 286 1543 294
rect 1483 269 1491 286
rect 1535 269 1543 286
rect 1483 250 1543 269
rect 1572 286 1632 294
rect 1572 269 1580 286
rect 1624 269 1632 286
rect 1572 250 1632 269
rect 1661 286 1721 294
rect 1661 269 1669 286
rect 1713 269 1721 286
rect 1661 250 1721 269
rect 1750 286 1810 294
rect 1750 269 1758 286
rect 1802 269 1810 286
rect 1750 250 1810 269
rect 1839 286 1899 294
rect 1839 269 1847 286
rect 1891 269 1899 286
rect 1839 250 1899 269
rect 1928 286 1988 294
rect 1928 269 1936 286
rect 1980 269 1988 286
rect 1928 250 1988 269
rect 2017 286 2077 294
rect 2017 269 2025 286
rect 2069 269 2077 286
rect 2017 250 2077 269
rect -2077 -269 -2017 -250
rect -2077 -286 -2069 -269
rect -2025 -286 -2017 -269
rect -2077 -294 -2017 -286
rect -1988 -269 -1928 -250
rect -1988 -286 -1980 -269
rect -1936 -286 -1928 -269
rect -1988 -294 -1928 -286
rect -1899 -269 -1839 -250
rect -1899 -286 -1891 -269
rect -1847 -286 -1839 -269
rect -1899 -294 -1839 -286
rect -1810 -269 -1750 -250
rect -1810 -286 -1802 -269
rect -1758 -286 -1750 -269
rect -1810 -294 -1750 -286
rect -1721 -269 -1661 -250
rect -1721 -286 -1713 -269
rect -1669 -286 -1661 -269
rect -1721 -294 -1661 -286
rect -1632 -269 -1572 -250
rect -1632 -286 -1624 -269
rect -1580 -286 -1572 -269
rect -1632 -294 -1572 -286
rect -1543 -269 -1483 -250
rect -1543 -286 -1535 -269
rect -1491 -286 -1483 -269
rect -1543 -294 -1483 -286
rect -1454 -269 -1394 -250
rect -1454 -286 -1446 -269
rect -1402 -286 -1394 -269
rect -1454 -294 -1394 -286
rect -1365 -269 -1305 -250
rect -1365 -286 -1357 -269
rect -1313 -286 -1305 -269
rect -1365 -294 -1305 -286
rect -1276 -269 -1216 -250
rect -1276 -286 -1268 -269
rect -1224 -286 -1216 -269
rect -1276 -294 -1216 -286
rect -1187 -269 -1127 -250
rect -1187 -286 -1179 -269
rect -1135 -286 -1127 -269
rect -1187 -294 -1127 -286
rect -1098 -269 -1038 -250
rect -1098 -286 -1090 -269
rect -1046 -286 -1038 -269
rect -1098 -294 -1038 -286
rect -1009 -269 -949 -250
rect -1009 -286 -1001 -269
rect -957 -286 -949 -269
rect -1009 -294 -949 -286
rect -920 -269 -860 -250
rect -920 -286 -912 -269
rect -868 -286 -860 -269
rect -920 -294 -860 -286
rect -831 -269 -771 -250
rect -831 -286 -823 -269
rect -779 -286 -771 -269
rect -831 -294 -771 -286
rect -742 -269 -682 -250
rect -742 -286 -734 -269
rect -690 -286 -682 -269
rect -742 -294 -682 -286
rect -653 -269 -593 -250
rect -653 -286 -645 -269
rect -601 -286 -593 -269
rect -653 -294 -593 -286
rect -564 -269 -504 -250
rect -564 -286 -556 -269
rect -512 -286 -504 -269
rect -564 -294 -504 -286
rect -475 -269 -415 -250
rect -475 -286 -467 -269
rect -423 -286 -415 -269
rect -475 -294 -415 -286
rect -386 -269 -326 -250
rect -386 -286 -378 -269
rect -334 -286 -326 -269
rect -386 -294 -326 -286
rect -297 -269 -237 -250
rect -297 -286 -289 -269
rect -245 -286 -237 -269
rect -297 -294 -237 -286
rect -208 -269 -148 -250
rect -208 -286 -200 -269
rect -156 -286 -148 -269
rect -208 -294 -148 -286
rect -119 -269 -59 -250
rect -119 -286 -111 -269
rect -67 -286 -59 -269
rect -119 -294 -59 -286
rect -30 -269 30 -250
rect -30 -286 -22 -269
rect 22 -286 30 -269
rect -30 -294 30 -286
rect 59 -269 119 -250
rect 59 -286 67 -269
rect 111 -286 119 -269
rect 59 -294 119 -286
rect 148 -269 208 -250
rect 148 -286 156 -269
rect 200 -286 208 -269
rect 148 -294 208 -286
rect 237 -269 297 -250
rect 237 -286 245 -269
rect 289 -286 297 -269
rect 237 -294 297 -286
rect 326 -269 386 -250
rect 326 -286 334 -269
rect 378 -286 386 -269
rect 326 -294 386 -286
rect 415 -269 475 -250
rect 415 -286 423 -269
rect 467 -286 475 -269
rect 415 -294 475 -286
rect 504 -269 564 -250
rect 504 -286 512 -269
rect 556 -286 564 -269
rect 504 -294 564 -286
rect 593 -269 653 -250
rect 593 -286 601 -269
rect 645 -286 653 -269
rect 593 -294 653 -286
rect 682 -269 742 -250
rect 682 -286 690 -269
rect 734 -286 742 -269
rect 682 -294 742 -286
rect 771 -269 831 -250
rect 771 -286 779 -269
rect 823 -286 831 -269
rect 771 -294 831 -286
rect 860 -269 920 -250
rect 860 -286 868 -269
rect 912 -286 920 -269
rect 860 -294 920 -286
rect 949 -269 1009 -250
rect 949 -286 957 -269
rect 1001 -286 1009 -269
rect 949 -294 1009 -286
rect 1038 -269 1098 -250
rect 1038 -286 1046 -269
rect 1090 -286 1098 -269
rect 1038 -294 1098 -286
rect 1127 -269 1187 -250
rect 1127 -286 1135 -269
rect 1179 -286 1187 -269
rect 1127 -294 1187 -286
rect 1216 -269 1276 -250
rect 1216 -286 1224 -269
rect 1268 -286 1276 -269
rect 1216 -294 1276 -286
rect 1305 -269 1365 -250
rect 1305 -286 1313 -269
rect 1357 -286 1365 -269
rect 1305 -294 1365 -286
rect 1394 -269 1454 -250
rect 1394 -286 1402 -269
rect 1446 -286 1454 -269
rect 1394 -294 1454 -286
rect 1483 -269 1543 -250
rect 1483 -286 1491 -269
rect 1535 -286 1543 -269
rect 1483 -294 1543 -286
rect 1572 -269 1632 -250
rect 1572 -286 1580 -269
rect 1624 -286 1632 -269
rect 1572 -294 1632 -286
rect 1661 -269 1721 -250
rect 1661 -286 1669 -269
rect 1713 -286 1721 -269
rect 1661 -294 1721 -286
rect 1750 -269 1810 -250
rect 1750 -286 1758 -269
rect 1802 -286 1810 -269
rect 1750 -294 1810 -286
rect 1839 -269 1899 -250
rect 1839 -286 1847 -269
rect 1891 -286 1899 -269
rect 1839 -294 1899 -286
rect 1928 -269 1988 -250
rect 1928 -286 1936 -269
rect 1980 -286 1988 -269
rect 1928 -294 1988 -286
rect 2017 -269 2077 -250
rect 2017 -286 2025 -269
rect 2069 -286 2077 -269
rect 2017 -294 2077 -286
<< polycont >>
rect -2069 269 -2025 286
rect -1980 269 -1936 286
rect -1891 269 -1847 286
rect -1802 269 -1758 286
rect -1713 269 -1669 286
rect -1624 269 -1580 286
rect -1535 269 -1491 286
rect -1446 269 -1402 286
rect -1357 269 -1313 286
rect -1268 269 -1224 286
rect -1179 269 -1135 286
rect -1090 269 -1046 286
rect -1001 269 -957 286
rect -912 269 -868 286
rect -823 269 -779 286
rect -734 269 -690 286
rect -645 269 -601 286
rect -556 269 -512 286
rect -467 269 -423 286
rect -378 269 -334 286
rect -289 269 -245 286
rect -200 269 -156 286
rect -111 269 -67 286
rect -22 269 22 286
rect 67 269 111 286
rect 156 269 200 286
rect 245 269 289 286
rect 334 269 378 286
rect 423 269 467 286
rect 512 269 556 286
rect 601 269 645 286
rect 690 269 734 286
rect 779 269 823 286
rect 868 269 912 286
rect 957 269 1001 286
rect 1046 269 1090 286
rect 1135 269 1179 286
rect 1224 269 1268 286
rect 1313 269 1357 286
rect 1402 269 1446 286
rect 1491 269 1535 286
rect 1580 269 1624 286
rect 1669 269 1713 286
rect 1758 269 1802 286
rect 1847 269 1891 286
rect 1936 269 1980 286
rect 2025 269 2069 286
rect -2069 -286 -2025 -269
rect -1980 -286 -1936 -269
rect -1891 -286 -1847 -269
rect -1802 -286 -1758 -269
rect -1713 -286 -1669 -269
rect -1624 -286 -1580 -269
rect -1535 -286 -1491 -269
rect -1446 -286 -1402 -269
rect -1357 -286 -1313 -269
rect -1268 -286 -1224 -269
rect -1179 -286 -1135 -269
rect -1090 -286 -1046 -269
rect -1001 -286 -957 -269
rect -912 -286 -868 -269
rect -823 -286 -779 -269
rect -734 -286 -690 -269
rect -645 -286 -601 -269
rect -556 -286 -512 -269
rect -467 -286 -423 -269
rect -378 -286 -334 -269
rect -289 -286 -245 -269
rect -200 -286 -156 -269
rect -111 -286 -67 -269
rect -22 -286 22 -269
rect 67 -286 111 -269
rect 156 -286 200 -269
rect 245 -286 289 -269
rect 334 -286 378 -269
rect 423 -286 467 -269
rect 512 -286 556 -269
rect 601 -286 645 -269
rect 690 -286 734 -269
rect 779 -286 823 -269
rect 868 -286 912 -269
rect 957 -286 1001 -269
rect 1046 -286 1090 -269
rect 1135 -286 1179 -269
rect 1224 -286 1268 -269
rect 1313 -286 1357 -269
rect 1402 -286 1446 -269
rect 1491 -286 1535 -269
rect 1580 -286 1624 -269
rect 1669 -286 1713 -269
rect 1758 -286 1802 -269
rect 1847 -286 1891 -269
rect 1936 -286 1980 -269
rect 2025 -286 2069 -269
<< locali >>
rect -2167 338 -2119 355
rect 2119 338 2167 355
rect -2167 307 -2150 338
rect 2150 307 2167 338
rect -2077 269 -2069 286
rect -2025 269 -2017 286
rect -1988 269 -1980 286
rect -1936 269 -1928 286
rect -1899 269 -1891 286
rect -1847 269 -1839 286
rect -1810 269 -1802 286
rect -1758 269 -1750 286
rect -1721 269 -1713 286
rect -1669 269 -1661 286
rect -1632 269 -1624 286
rect -1580 269 -1572 286
rect -1543 269 -1535 286
rect -1491 269 -1483 286
rect -1454 269 -1446 286
rect -1402 269 -1394 286
rect -1365 269 -1357 286
rect -1313 269 -1305 286
rect -1276 269 -1268 286
rect -1224 269 -1216 286
rect -1187 269 -1179 286
rect -1135 269 -1127 286
rect -1098 269 -1090 286
rect -1046 269 -1038 286
rect -1009 269 -1001 286
rect -957 269 -949 286
rect -920 269 -912 286
rect -868 269 -860 286
rect -831 269 -823 286
rect -779 269 -771 286
rect -742 269 -734 286
rect -690 269 -682 286
rect -653 269 -645 286
rect -601 269 -593 286
rect -564 269 -556 286
rect -512 269 -504 286
rect -475 269 -467 286
rect -423 269 -415 286
rect -386 269 -378 286
rect -334 269 -326 286
rect -297 269 -289 286
rect -245 269 -237 286
rect -208 269 -200 286
rect -156 269 -148 286
rect -119 269 -111 286
rect -67 269 -59 286
rect -30 269 -22 286
rect 22 269 30 286
rect 59 269 67 286
rect 111 269 119 286
rect 148 269 156 286
rect 200 269 208 286
rect 237 269 245 286
rect 289 269 297 286
rect 326 269 334 286
rect 378 269 386 286
rect 415 269 423 286
rect 467 269 475 286
rect 504 269 512 286
rect 556 269 564 286
rect 593 269 601 286
rect 645 269 653 286
rect 682 269 690 286
rect 734 269 742 286
rect 771 269 779 286
rect 823 269 831 286
rect 860 269 868 286
rect 912 269 920 286
rect 949 269 957 286
rect 1001 269 1009 286
rect 1038 269 1046 286
rect 1090 269 1098 286
rect 1127 269 1135 286
rect 1179 269 1187 286
rect 1216 269 1224 286
rect 1268 269 1276 286
rect 1305 269 1313 286
rect 1357 269 1365 286
rect 1394 269 1402 286
rect 1446 269 1454 286
rect 1483 269 1491 286
rect 1535 269 1543 286
rect 1572 269 1580 286
rect 1624 269 1632 286
rect 1661 269 1669 286
rect 1713 269 1721 286
rect 1750 269 1758 286
rect 1802 269 1810 286
rect 1839 269 1847 286
rect 1891 269 1899 286
rect 1928 269 1936 286
rect 1980 269 1988 286
rect 2017 269 2025 286
rect 2069 269 2077 286
rect -2100 244 -2083 252
rect -2100 -252 -2083 -244
rect -2011 244 -1994 252
rect -2011 -252 -1994 -244
rect -1922 244 -1905 252
rect -1922 -252 -1905 -244
rect -1833 244 -1816 252
rect -1833 -252 -1816 -244
rect -1744 244 -1727 252
rect -1744 -252 -1727 -244
rect -1655 244 -1638 252
rect -1655 -252 -1638 -244
rect -1566 244 -1549 252
rect -1566 -252 -1549 -244
rect -1477 244 -1460 252
rect -1477 -252 -1460 -244
rect -1388 244 -1371 252
rect -1388 -252 -1371 -244
rect -1299 244 -1282 252
rect -1299 -252 -1282 -244
rect -1210 244 -1193 252
rect -1210 -252 -1193 -244
rect -1121 244 -1104 252
rect -1121 -252 -1104 -244
rect -1032 244 -1015 252
rect -1032 -252 -1015 -244
rect -943 244 -926 252
rect -943 -252 -926 -244
rect -854 244 -837 252
rect -854 -252 -837 -244
rect -765 244 -748 252
rect -765 -252 -748 -244
rect -676 244 -659 252
rect -676 -252 -659 -244
rect -587 244 -570 252
rect -587 -252 -570 -244
rect -498 244 -481 252
rect -498 -252 -481 -244
rect -409 244 -392 252
rect -409 -252 -392 -244
rect -320 244 -303 252
rect -320 -252 -303 -244
rect -231 244 -214 252
rect -231 -252 -214 -244
rect -142 244 -125 252
rect -142 -252 -125 -244
rect -53 244 -36 252
rect -53 -252 -36 -244
rect 36 244 53 252
rect 36 -252 53 -244
rect 125 244 142 252
rect 125 -252 142 -244
rect 214 244 231 252
rect 214 -252 231 -244
rect 303 244 320 252
rect 303 -252 320 -244
rect 392 244 409 252
rect 392 -252 409 -244
rect 481 244 498 252
rect 481 -252 498 -244
rect 570 244 587 252
rect 570 -252 587 -244
rect 659 244 676 252
rect 659 -252 676 -244
rect 748 244 765 252
rect 748 -252 765 -244
rect 837 244 854 252
rect 837 -252 854 -244
rect 926 244 943 252
rect 926 -252 943 -244
rect 1015 244 1032 252
rect 1015 -252 1032 -244
rect 1104 244 1121 252
rect 1104 -252 1121 -244
rect 1193 244 1210 252
rect 1193 -252 1210 -244
rect 1282 244 1299 252
rect 1282 -252 1299 -244
rect 1371 244 1388 252
rect 1371 -252 1388 -244
rect 1460 244 1477 252
rect 1460 -252 1477 -244
rect 1549 244 1566 252
rect 1549 -252 1566 -244
rect 1638 244 1655 252
rect 1638 -252 1655 -244
rect 1727 244 1744 252
rect 1727 -252 1744 -244
rect 1816 244 1833 252
rect 1816 -252 1833 -244
rect 1905 244 1922 252
rect 1905 -252 1922 -244
rect 1994 244 2011 252
rect 1994 -252 2011 -244
rect 2083 244 2100 252
rect 2083 -252 2100 -244
rect -2077 -286 -2069 -269
rect -2025 -286 -2017 -269
rect -1988 -286 -1980 -269
rect -1936 -286 -1928 -269
rect -1899 -286 -1891 -269
rect -1847 -286 -1839 -269
rect -1810 -286 -1802 -269
rect -1758 -286 -1750 -269
rect -1721 -286 -1713 -269
rect -1669 -286 -1661 -269
rect -1632 -286 -1624 -269
rect -1580 -286 -1572 -269
rect -1543 -286 -1535 -269
rect -1491 -286 -1483 -269
rect -1454 -286 -1446 -269
rect -1402 -286 -1394 -269
rect -1365 -286 -1357 -269
rect -1313 -286 -1305 -269
rect -1276 -286 -1268 -269
rect -1224 -286 -1216 -269
rect -1187 -286 -1179 -269
rect -1135 -286 -1127 -269
rect -1098 -286 -1090 -269
rect -1046 -286 -1038 -269
rect -1009 -286 -1001 -269
rect -957 -286 -949 -269
rect -920 -286 -912 -269
rect -868 -286 -860 -269
rect -831 -286 -823 -269
rect -779 -286 -771 -269
rect -742 -286 -734 -269
rect -690 -286 -682 -269
rect -653 -286 -645 -269
rect -601 -286 -593 -269
rect -564 -286 -556 -269
rect -512 -286 -504 -269
rect -475 -286 -467 -269
rect -423 -286 -415 -269
rect -386 -286 -378 -269
rect -334 -286 -326 -269
rect -297 -286 -289 -269
rect -245 -286 -237 -269
rect -208 -286 -200 -269
rect -156 -286 -148 -269
rect -119 -286 -111 -269
rect -67 -286 -59 -269
rect -30 -286 -22 -269
rect 22 -286 30 -269
rect 59 -286 67 -269
rect 111 -286 119 -269
rect 148 -286 156 -269
rect 200 -286 208 -269
rect 237 -286 245 -269
rect 289 -286 297 -269
rect 326 -286 334 -269
rect 378 -286 386 -269
rect 415 -286 423 -269
rect 467 -286 475 -269
rect 504 -286 512 -269
rect 556 -286 564 -269
rect 593 -286 601 -269
rect 645 -286 653 -269
rect 682 -286 690 -269
rect 734 -286 742 -269
rect 771 -286 779 -269
rect 823 -286 831 -269
rect 860 -286 868 -269
rect 912 -286 920 -269
rect 949 -286 957 -269
rect 1001 -286 1009 -269
rect 1038 -286 1046 -269
rect 1090 -286 1098 -269
rect 1127 -286 1135 -269
rect 1179 -286 1187 -269
rect 1216 -286 1224 -269
rect 1268 -286 1276 -269
rect 1305 -286 1313 -269
rect 1357 -286 1365 -269
rect 1394 -286 1402 -269
rect 1446 -286 1454 -269
rect 1483 -286 1491 -269
rect 1535 -286 1543 -269
rect 1572 -286 1580 -269
rect 1624 -286 1632 -269
rect 1661 -286 1669 -269
rect 1713 -286 1721 -269
rect 1750 -286 1758 -269
rect 1802 -286 1810 -269
rect 1839 -286 1847 -269
rect 1891 -286 1899 -269
rect 1928 -286 1936 -269
rect 1980 -286 1988 -269
rect 2017 -286 2025 -269
rect 2069 -286 2077 -269
rect -2167 -338 -2150 -307
rect 2150 -338 2167 -307
rect -2167 -355 -2119 -338
rect 2119 -355 2167 -338
<< viali >>
rect -2069 269 -2025 286
rect -1980 269 -1936 286
rect -1891 269 -1847 286
rect -1802 269 -1758 286
rect -1713 269 -1669 286
rect -1624 269 -1580 286
rect -1535 269 -1491 286
rect -1446 269 -1402 286
rect -1357 269 -1313 286
rect -1268 269 -1224 286
rect -1179 269 -1135 286
rect -1090 269 -1046 286
rect -1001 269 -957 286
rect -912 269 -868 286
rect -823 269 -779 286
rect -734 269 -690 286
rect -645 269 -601 286
rect -556 269 -512 286
rect -467 269 -423 286
rect -378 269 -334 286
rect -289 269 -245 286
rect -200 269 -156 286
rect -111 269 -67 286
rect -22 269 22 286
rect 67 269 111 286
rect 156 269 200 286
rect 245 269 289 286
rect 334 269 378 286
rect 423 269 467 286
rect 512 269 556 286
rect 601 269 645 286
rect 690 269 734 286
rect 779 269 823 286
rect 868 269 912 286
rect 957 269 1001 286
rect 1046 269 1090 286
rect 1135 269 1179 286
rect 1224 269 1268 286
rect 1313 269 1357 286
rect 1402 269 1446 286
rect 1491 269 1535 286
rect 1580 269 1624 286
rect 1669 269 1713 286
rect 1758 269 1802 286
rect 1847 269 1891 286
rect 1936 269 1980 286
rect 2025 269 2069 286
rect -2100 -244 -2083 244
rect -2011 -244 -1994 244
rect -1922 -244 -1905 244
rect -1833 -244 -1816 244
rect -1744 -244 -1727 244
rect -1655 -244 -1638 244
rect -1566 -244 -1549 244
rect -1477 -244 -1460 244
rect -1388 -244 -1371 244
rect -1299 -244 -1282 244
rect -1210 -244 -1193 244
rect -1121 -244 -1104 244
rect -1032 -244 -1015 244
rect -943 -244 -926 244
rect -854 -244 -837 244
rect -765 -244 -748 244
rect -676 -244 -659 244
rect -587 -244 -570 244
rect -498 -244 -481 244
rect -409 -244 -392 244
rect -320 -244 -303 244
rect -231 -244 -214 244
rect -142 -244 -125 244
rect -53 -244 -36 244
rect 36 -244 53 244
rect 125 -244 142 244
rect 214 -244 231 244
rect 303 -244 320 244
rect 392 -244 409 244
rect 481 -244 498 244
rect 570 -244 587 244
rect 659 -244 676 244
rect 748 -244 765 244
rect 837 -244 854 244
rect 926 -244 943 244
rect 1015 -244 1032 244
rect 1104 -244 1121 244
rect 1193 -244 1210 244
rect 1282 -244 1299 244
rect 1371 -244 1388 244
rect 1460 -244 1477 244
rect 1549 -244 1566 244
rect 1638 -244 1655 244
rect 1727 -244 1744 244
rect 1816 -244 1833 244
rect 1905 -244 1922 244
rect 1994 -244 2011 244
rect 2083 -244 2100 244
rect -2069 -286 -2025 -269
rect -1980 -286 -1936 -269
rect -1891 -286 -1847 -269
rect -1802 -286 -1758 -269
rect -1713 -286 -1669 -269
rect -1624 -286 -1580 -269
rect -1535 -286 -1491 -269
rect -1446 -286 -1402 -269
rect -1357 -286 -1313 -269
rect -1268 -286 -1224 -269
rect -1179 -286 -1135 -269
rect -1090 -286 -1046 -269
rect -1001 -286 -957 -269
rect -912 -286 -868 -269
rect -823 -286 -779 -269
rect -734 -286 -690 -269
rect -645 -286 -601 -269
rect -556 -286 -512 -269
rect -467 -286 -423 -269
rect -378 -286 -334 -269
rect -289 -286 -245 -269
rect -200 -286 -156 -269
rect -111 -286 -67 -269
rect -22 -286 22 -269
rect 67 -286 111 -269
rect 156 -286 200 -269
rect 245 -286 289 -269
rect 334 -286 378 -269
rect 423 -286 467 -269
rect 512 -286 556 -269
rect 601 -286 645 -269
rect 690 -286 734 -269
rect 779 -286 823 -269
rect 868 -286 912 -269
rect 957 -286 1001 -269
rect 1046 -286 1090 -269
rect 1135 -286 1179 -269
rect 1224 -286 1268 -269
rect 1313 -286 1357 -269
rect 1402 -286 1446 -269
rect 1491 -286 1535 -269
rect 1580 -286 1624 -269
rect 1669 -286 1713 -269
rect 1758 -286 1802 -269
rect 1847 -286 1891 -269
rect 1936 -286 1980 -269
rect 2025 -286 2069 -269
<< metal1 >>
rect -2075 286 -2019 289
rect -2075 269 -2069 286
rect -2025 269 -2019 286
rect -2075 266 -2019 269
rect -1986 286 -1930 289
rect -1986 269 -1980 286
rect -1936 269 -1930 286
rect -1986 266 -1930 269
rect -1897 286 -1841 289
rect -1897 269 -1891 286
rect -1847 269 -1841 286
rect -1897 266 -1841 269
rect -1808 286 -1752 289
rect -1808 269 -1802 286
rect -1758 269 -1752 286
rect -1808 266 -1752 269
rect -1719 286 -1663 289
rect -1719 269 -1713 286
rect -1669 269 -1663 286
rect -1719 266 -1663 269
rect -1630 286 -1574 289
rect -1630 269 -1624 286
rect -1580 269 -1574 286
rect -1630 266 -1574 269
rect -1541 286 -1485 289
rect -1541 269 -1535 286
rect -1491 269 -1485 286
rect -1541 266 -1485 269
rect -1452 286 -1396 289
rect -1452 269 -1446 286
rect -1402 269 -1396 286
rect -1452 266 -1396 269
rect -1363 286 -1307 289
rect -1363 269 -1357 286
rect -1313 269 -1307 286
rect -1363 266 -1307 269
rect -1274 286 -1218 289
rect -1274 269 -1268 286
rect -1224 269 -1218 286
rect -1274 266 -1218 269
rect -1185 286 -1129 289
rect -1185 269 -1179 286
rect -1135 269 -1129 286
rect -1185 266 -1129 269
rect -1096 286 -1040 289
rect -1096 269 -1090 286
rect -1046 269 -1040 286
rect -1096 266 -1040 269
rect -1007 286 -951 289
rect -1007 269 -1001 286
rect -957 269 -951 286
rect -1007 266 -951 269
rect -918 286 -862 289
rect -918 269 -912 286
rect -868 269 -862 286
rect -918 266 -862 269
rect -829 286 -773 289
rect -829 269 -823 286
rect -779 269 -773 286
rect -829 266 -773 269
rect -740 286 -684 289
rect -740 269 -734 286
rect -690 269 -684 286
rect -740 266 -684 269
rect -651 286 -595 289
rect -651 269 -645 286
rect -601 269 -595 286
rect -651 266 -595 269
rect -562 286 -506 289
rect -562 269 -556 286
rect -512 269 -506 286
rect -562 266 -506 269
rect -473 286 -417 289
rect -473 269 -467 286
rect -423 269 -417 286
rect -473 266 -417 269
rect -384 286 -328 289
rect -384 269 -378 286
rect -334 269 -328 286
rect -384 266 -328 269
rect -295 286 -239 289
rect -295 269 -289 286
rect -245 269 -239 286
rect -295 266 -239 269
rect -206 286 -150 289
rect -206 269 -200 286
rect -156 269 -150 286
rect -206 266 -150 269
rect -117 286 -61 289
rect -117 269 -111 286
rect -67 269 -61 286
rect -117 266 -61 269
rect -28 286 28 289
rect -28 269 -22 286
rect 22 269 28 286
rect -28 266 28 269
rect 61 286 117 289
rect 61 269 67 286
rect 111 269 117 286
rect 61 266 117 269
rect 150 286 206 289
rect 150 269 156 286
rect 200 269 206 286
rect 150 266 206 269
rect 239 286 295 289
rect 239 269 245 286
rect 289 269 295 286
rect 239 266 295 269
rect 328 286 384 289
rect 328 269 334 286
rect 378 269 384 286
rect 328 266 384 269
rect 417 286 473 289
rect 417 269 423 286
rect 467 269 473 286
rect 417 266 473 269
rect 506 286 562 289
rect 506 269 512 286
rect 556 269 562 286
rect 506 266 562 269
rect 595 286 651 289
rect 595 269 601 286
rect 645 269 651 286
rect 595 266 651 269
rect 684 286 740 289
rect 684 269 690 286
rect 734 269 740 286
rect 684 266 740 269
rect 773 286 829 289
rect 773 269 779 286
rect 823 269 829 286
rect 773 266 829 269
rect 862 286 918 289
rect 862 269 868 286
rect 912 269 918 286
rect 862 266 918 269
rect 951 286 1007 289
rect 951 269 957 286
rect 1001 269 1007 286
rect 951 266 1007 269
rect 1040 286 1096 289
rect 1040 269 1046 286
rect 1090 269 1096 286
rect 1040 266 1096 269
rect 1129 286 1185 289
rect 1129 269 1135 286
rect 1179 269 1185 286
rect 1129 266 1185 269
rect 1218 286 1274 289
rect 1218 269 1224 286
rect 1268 269 1274 286
rect 1218 266 1274 269
rect 1307 286 1363 289
rect 1307 269 1313 286
rect 1357 269 1363 286
rect 1307 266 1363 269
rect 1396 286 1452 289
rect 1396 269 1402 286
rect 1446 269 1452 286
rect 1396 266 1452 269
rect 1485 286 1541 289
rect 1485 269 1491 286
rect 1535 269 1541 286
rect 1485 266 1541 269
rect 1574 286 1630 289
rect 1574 269 1580 286
rect 1624 269 1630 286
rect 1574 266 1630 269
rect 1663 286 1719 289
rect 1663 269 1669 286
rect 1713 269 1719 286
rect 1663 266 1719 269
rect 1752 286 1808 289
rect 1752 269 1758 286
rect 1802 269 1808 286
rect 1752 266 1808 269
rect 1841 286 1897 289
rect 1841 269 1847 286
rect 1891 269 1897 286
rect 1841 266 1897 269
rect 1930 286 1986 289
rect 1930 269 1936 286
rect 1980 269 1986 286
rect 1930 266 1986 269
rect 2019 286 2075 289
rect 2019 269 2025 286
rect 2069 269 2075 286
rect 2019 266 2075 269
rect -2103 244 -2080 250
rect -2103 -244 -2100 244
rect -2083 -244 -2080 244
rect -2103 -250 -2080 -244
rect -2014 244 -1991 250
rect -2014 -244 -2011 244
rect -1994 -244 -1991 244
rect -2014 -250 -1991 -244
rect -1925 244 -1902 250
rect -1925 -244 -1922 244
rect -1905 -244 -1902 244
rect -1925 -250 -1902 -244
rect -1836 244 -1813 250
rect -1836 -244 -1833 244
rect -1816 -244 -1813 244
rect -1836 -250 -1813 -244
rect -1747 244 -1724 250
rect -1747 -244 -1744 244
rect -1727 -244 -1724 244
rect -1747 -250 -1724 -244
rect -1658 244 -1635 250
rect -1658 -244 -1655 244
rect -1638 -244 -1635 244
rect -1658 -250 -1635 -244
rect -1569 244 -1546 250
rect -1569 -244 -1566 244
rect -1549 -244 -1546 244
rect -1569 -250 -1546 -244
rect -1480 244 -1457 250
rect -1480 -244 -1477 244
rect -1460 -244 -1457 244
rect -1480 -250 -1457 -244
rect -1391 244 -1368 250
rect -1391 -244 -1388 244
rect -1371 -244 -1368 244
rect -1391 -250 -1368 -244
rect -1302 244 -1279 250
rect -1302 -244 -1299 244
rect -1282 -244 -1279 244
rect -1302 -250 -1279 -244
rect -1213 244 -1190 250
rect -1213 -244 -1210 244
rect -1193 -244 -1190 244
rect -1213 -250 -1190 -244
rect -1124 244 -1101 250
rect -1124 -244 -1121 244
rect -1104 -244 -1101 244
rect -1124 -250 -1101 -244
rect -1035 244 -1012 250
rect -1035 -244 -1032 244
rect -1015 -244 -1012 244
rect -1035 -250 -1012 -244
rect -946 244 -923 250
rect -946 -244 -943 244
rect -926 -244 -923 244
rect -946 -250 -923 -244
rect -857 244 -834 250
rect -857 -244 -854 244
rect -837 -244 -834 244
rect -857 -250 -834 -244
rect -768 244 -745 250
rect -768 -244 -765 244
rect -748 -244 -745 244
rect -768 -250 -745 -244
rect -679 244 -656 250
rect -679 -244 -676 244
rect -659 -244 -656 244
rect -679 -250 -656 -244
rect -590 244 -567 250
rect -590 -244 -587 244
rect -570 -244 -567 244
rect -590 -250 -567 -244
rect -501 244 -478 250
rect -501 -244 -498 244
rect -481 -244 -478 244
rect -501 -250 -478 -244
rect -412 244 -389 250
rect -412 -244 -409 244
rect -392 -244 -389 244
rect -412 -250 -389 -244
rect -323 244 -300 250
rect -323 -244 -320 244
rect -303 -244 -300 244
rect -323 -250 -300 -244
rect -234 244 -211 250
rect -234 -244 -231 244
rect -214 -244 -211 244
rect -234 -250 -211 -244
rect -145 244 -122 250
rect -145 -244 -142 244
rect -125 -244 -122 244
rect -145 -250 -122 -244
rect -56 244 -33 250
rect -56 -244 -53 244
rect -36 -244 -33 244
rect -56 -250 -33 -244
rect 33 244 56 250
rect 33 -244 36 244
rect 53 -244 56 244
rect 33 -250 56 -244
rect 122 244 145 250
rect 122 -244 125 244
rect 142 -244 145 244
rect 122 -250 145 -244
rect 211 244 234 250
rect 211 -244 214 244
rect 231 -244 234 244
rect 211 -250 234 -244
rect 300 244 323 250
rect 300 -244 303 244
rect 320 -244 323 244
rect 300 -250 323 -244
rect 389 244 412 250
rect 389 -244 392 244
rect 409 -244 412 244
rect 389 -250 412 -244
rect 478 244 501 250
rect 478 -244 481 244
rect 498 -244 501 244
rect 478 -250 501 -244
rect 567 244 590 250
rect 567 -244 570 244
rect 587 -244 590 244
rect 567 -250 590 -244
rect 656 244 679 250
rect 656 -244 659 244
rect 676 -244 679 244
rect 656 -250 679 -244
rect 745 244 768 250
rect 745 -244 748 244
rect 765 -244 768 244
rect 745 -250 768 -244
rect 834 244 857 250
rect 834 -244 837 244
rect 854 -244 857 244
rect 834 -250 857 -244
rect 923 244 946 250
rect 923 -244 926 244
rect 943 -244 946 244
rect 923 -250 946 -244
rect 1012 244 1035 250
rect 1012 -244 1015 244
rect 1032 -244 1035 244
rect 1012 -250 1035 -244
rect 1101 244 1124 250
rect 1101 -244 1104 244
rect 1121 -244 1124 244
rect 1101 -250 1124 -244
rect 1190 244 1213 250
rect 1190 -244 1193 244
rect 1210 -244 1213 244
rect 1190 -250 1213 -244
rect 1279 244 1302 250
rect 1279 -244 1282 244
rect 1299 -244 1302 244
rect 1279 -250 1302 -244
rect 1368 244 1391 250
rect 1368 -244 1371 244
rect 1388 -244 1391 244
rect 1368 -250 1391 -244
rect 1457 244 1480 250
rect 1457 -244 1460 244
rect 1477 -244 1480 244
rect 1457 -250 1480 -244
rect 1546 244 1569 250
rect 1546 -244 1549 244
rect 1566 -244 1569 244
rect 1546 -250 1569 -244
rect 1635 244 1658 250
rect 1635 -244 1638 244
rect 1655 -244 1658 244
rect 1635 -250 1658 -244
rect 1724 244 1747 250
rect 1724 -244 1727 244
rect 1744 -244 1747 244
rect 1724 -250 1747 -244
rect 1813 244 1836 250
rect 1813 -244 1816 244
rect 1833 -244 1836 244
rect 1813 -250 1836 -244
rect 1902 244 1925 250
rect 1902 -244 1905 244
rect 1922 -244 1925 244
rect 1902 -250 1925 -244
rect 1991 244 2014 250
rect 1991 -244 1994 244
rect 2011 -244 2014 244
rect 1991 -250 2014 -244
rect 2080 244 2103 250
rect 2080 -244 2083 244
rect 2100 -244 2103 244
rect 2080 -250 2103 -244
rect -2075 -269 -2019 -266
rect -2075 -286 -2069 -269
rect -2025 -286 -2019 -269
rect -2075 -289 -2019 -286
rect -1986 -269 -1930 -266
rect -1986 -286 -1980 -269
rect -1936 -286 -1930 -269
rect -1986 -289 -1930 -286
rect -1897 -269 -1841 -266
rect -1897 -286 -1891 -269
rect -1847 -286 -1841 -269
rect -1897 -289 -1841 -286
rect -1808 -269 -1752 -266
rect -1808 -286 -1802 -269
rect -1758 -286 -1752 -269
rect -1808 -289 -1752 -286
rect -1719 -269 -1663 -266
rect -1719 -286 -1713 -269
rect -1669 -286 -1663 -269
rect -1719 -289 -1663 -286
rect -1630 -269 -1574 -266
rect -1630 -286 -1624 -269
rect -1580 -286 -1574 -269
rect -1630 -289 -1574 -286
rect -1541 -269 -1485 -266
rect -1541 -286 -1535 -269
rect -1491 -286 -1485 -269
rect -1541 -289 -1485 -286
rect -1452 -269 -1396 -266
rect -1452 -286 -1446 -269
rect -1402 -286 -1396 -269
rect -1452 -289 -1396 -286
rect -1363 -269 -1307 -266
rect -1363 -286 -1357 -269
rect -1313 -286 -1307 -269
rect -1363 -289 -1307 -286
rect -1274 -269 -1218 -266
rect -1274 -286 -1268 -269
rect -1224 -286 -1218 -269
rect -1274 -289 -1218 -286
rect -1185 -269 -1129 -266
rect -1185 -286 -1179 -269
rect -1135 -286 -1129 -269
rect -1185 -289 -1129 -286
rect -1096 -269 -1040 -266
rect -1096 -286 -1090 -269
rect -1046 -286 -1040 -269
rect -1096 -289 -1040 -286
rect -1007 -269 -951 -266
rect -1007 -286 -1001 -269
rect -957 -286 -951 -269
rect -1007 -289 -951 -286
rect -918 -269 -862 -266
rect -918 -286 -912 -269
rect -868 -286 -862 -269
rect -918 -289 -862 -286
rect -829 -269 -773 -266
rect -829 -286 -823 -269
rect -779 -286 -773 -269
rect -829 -289 -773 -286
rect -740 -269 -684 -266
rect -740 -286 -734 -269
rect -690 -286 -684 -269
rect -740 -289 -684 -286
rect -651 -269 -595 -266
rect -651 -286 -645 -269
rect -601 -286 -595 -269
rect -651 -289 -595 -286
rect -562 -269 -506 -266
rect -562 -286 -556 -269
rect -512 -286 -506 -269
rect -562 -289 -506 -286
rect -473 -269 -417 -266
rect -473 -286 -467 -269
rect -423 -286 -417 -269
rect -473 -289 -417 -286
rect -384 -269 -328 -266
rect -384 -286 -378 -269
rect -334 -286 -328 -269
rect -384 -289 -328 -286
rect -295 -269 -239 -266
rect -295 -286 -289 -269
rect -245 -286 -239 -269
rect -295 -289 -239 -286
rect -206 -269 -150 -266
rect -206 -286 -200 -269
rect -156 -286 -150 -269
rect -206 -289 -150 -286
rect -117 -269 -61 -266
rect -117 -286 -111 -269
rect -67 -286 -61 -269
rect -117 -289 -61 -286
rect -28 -269 28 -266
rect -28 -286 -22 -269
rect 22 -286 28 -269
rect -28 -289 28 -286
rect 61 -269 117 -266
rect 61 -286 67 -269
rect 111 -286 117 -269
rect 61 -289 117 -286
rect 150 -269 206 -266
rect 150 -286 156 -269
rect 200 -286 206 -269
rect 150 -289 206 -286
rect 239 -269 295 -266
rect 239 -286 245 -269
rect 289 -286 295 -269
rect 239 -289 295 -286
rect 328 -269 384 -266
rect 328 -286 334 -269
rect 378 -286 384 -269
rect 328 -289 384 -286
rect 417 -269 473 -266
rect 417 -286 423 -269
rect 467 -286 473 -269
rect 417 -289 473 -286
rect 506 -269 562 -266
rect 506 -286 512 -269
rect 556 -286 562 -269
rect 506 -289 562 -286
rect 595 -269 651 -266
rect 595 -286 601 -269
rect 645 -286 651 -269
rect 595 -289 651 -286
rect 684 -269 740 -266
rect 684 -286 690 -269
rect 734 -286 740 -269
rect 684 -289 740 -286
rect 773 -269 829 -266
rect 773 -286 779 -269
rect 823 -286 829 -269
rect 773 -289 829 -286
rect 862 -269 918 -266
rect 862 -286 868 -269
rect 912 -286 918 -269
rect 862 -289 918 -286
rect 951 -269 1007 -266
rect 951 -286 957 -269
rect 1001 -286 1007 -269
rect 951 -289 1007 -286
rect 1040 -269 1096 -266
rect 1040 -286 1046 -269
rect 1090 -286 1096 -269
rect 1040 -289 1096 -286
rect 1129 -269 1185 -266
rect 1129 -286 1135 -269
rect 1179 -286 1185 -269
rect 1129 -289 1185 -286
rect 1218 -269 1274 -266
rect 1218 -286 1224 -269
rect 1268 -286 1274 -269
rect 1218 -289 1274 -286
rect 1307 -269 1363 -266
rect 1307 -286 1313 -269
rect 1357 -286 1363 -269
rect 1307 -289 1363 -286
rect 1396 -269 1452 -266
rect 1396 -286 1402 -269
rect 1446 -286 1452 -269
rect 1396 -289 1452 -286
rect 1485 -269 1541 -266
rect 1485 -286 1491 -269
rect 1535 -286 1541 -269
rect 1485 -289 1541 -286
rect 1574 -269 1630 -266
rect 1574 -286 1580 -269
rect 1624 -286 1630 -269
rect 1574 -289 1630 -286
rect 1663 -269 1719 -266
rect 1663 -286 1669 -269
rect 1713 -286 1719 -269
rect 1663 -289 1719 -286
rect 1752 -269 1808 -266
rect 1752 -286 1758 -269
rect 1802 -286 1808 -269
rect 1752 -289 1808 -286
rect 1841 -269 1897 -266
rect 1841 -286 1847 -269
rect 1891 -286 1897 -269
rect 1841 -289 1897 -286
rect 1930 -269 1986 -266
rect 1930 -286 1936 -269
rect 1980 -286 1986 -269
rect 1930 -289 1986 -286
rect 2019 -269 2075 -266
rect 2019 -286 2025 -269
rect 2069 -286 2075 -269
rect 2019 -289 2075 -286
<< properties >>
string FIXED_BBOX -2158 -346 2158 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.6 m 1 nf 47 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
