magic
tech sky130A
magscale 1 2
timestamp 1712014955
<< pwell >>
rect -1089 -327 1089 327
<< mvnmos >>
rect -861 -131 -741 69
rect -683 -131 -563 69
rect -505 -131 -385 69
rect -327 -131 -207 69
rect -149 -131 -29 69
rect 29 -131 149 69
rect 207 -131 327 69
rect 385 -131 505 69
rect 563 -131 683 69
rect 741 -131 861 69
<< mvndiff >>
rect -919 57 -861 69
rect -919 -119 -907 57
rect -873 -119 -861 57
rect -919 -131 -861 -119
rect -741 57 -683 69
rect -741 -119 -729 57
rect -695 -119 -683 57
rect -741 -131 -683 -119
rect -563 57 -505 69
rect -563 -119 -551 57
rect -517 -119 -505 57
rect -563 -131 -505 -119
rect -385 57 -327 69
rect -385 -119 -373 57
rect -339 -119 -327 57
rect -385 -131 -327 -119
rect -207 57 -149 69
rect -207 -119 -195 57
rect -161 -119 -149 57
rect -207 -131 -149 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 149 57 207 69
rect 149 -119 161 57
rect 195 -119 207 57
rect 149 -131 207 -119
rect 327 57 385 69
rect 327 -119 339 57
rect 373 -119 385 57
rect 327 -131 385 -119
rect 505 57 563 69
rect 505 -119 517 57
rect 551 -119 563 57
rect 505 -131 563 -119
rect 683 57 741 69
rect 683 -119 695 57
rect 729 -119 741 57
rect 683 -131 741 -119
rect 861 57 919 69
rect 861 -119 873 57
rect 907 -119 919 57
rect 861 -131 919 -119
<< mvndiffc >>
rect -907 -119 -873 57
rect -729 -119 -695 57
rect -551 -119 -517 57
rect -373 -119 -339 57
rect -195 -119 -161 57
rect -17 -119 17 57
rect 161 -119 195 57
rect 339 -119 373 57
rect 517 -119 551 57
rect 695 -119 729 57
rect 873 -119 907 57
<< mvpsubdiff >>
rect -1053 279 1053 291
rect -1053 245 -945 279
rect 945 245 1053 279
rect -1053 233 1053 245
rect -1053 183 -995 233
rect -1053 -183 -1041 183
rect -1007 -183 -995 183
rect 995 183 1053 233
rect -1053 -233 -995 -183
rect 995 -183 1007 183
rect 1041 -183 1053 183
rect 995 -233 1053 -183
rect -1053 -245 1053 -233
rect -1053 -279 -945 -245
rect 945 -279 1053 -245
rect -1053 -291 1053 -279
<< mvpsubdiffcont >>
rect -945 245 945 279
rect -1041 -183 -1007 183
rect 1007 -183 1041 183
rect -945 -279 945 -245
<< poly >>
rect -861 141 -741 157
rect -861 107 -845 141
rect -757 107 -741 141
rect -861 69 -741 107
rect -683 141 -563 157
rect -683 107 -667 141
rect -579 107 -563 141
rect -683 69 -563 107
rect -505 141 -385 157
rect -505 107 -489 141
rect -401 107 -385 141
rect -505 69 -385 107
rect -327 141 -207 157
rect -327 107 -311 141
rect -223 107 -207 141
rect -327 69 -207 107
rect -149 141 -29 157
rect -149 107 -133 141
rect -45 107 -29 141
rect -149 69 -29 107
rect 29 141 149 157
rect 29 107 45 141
rect 133 107 149 141
rect 29 69 149 107
rect 207 141 327 157
rect 207 107 223 141
rect 311 107 327 141
rect 207 69 327 107
rect 385 141 505 157
rect 385 107 401 141
rect 489 107 505 141
rect 385 69 505 107
rect 563 141 683 157
rect 563 107 579 141
rect 667 107 683 141
rect 563 69 683 107
rect 741 141 861 157
rect 741 107 757 141
rect 845 107 861 141
rect 741 69 861 107
rect -861 -157 -741 -131
rect -683 -157 -563 -131
rect -505 -157 -385 -131
rect -327 -157 -207 -131
rect -149 -157 -29 -131
rect 29 -157 149 -131
rect 207 -157 327 -131
rect 385 -157 505 -131
rect 563 -157 683 -131
rect 741 -157 861 -131
<< polycont >>
rect -845 107 -757 141
rect -667 107 -579 141
rect -489 107 -401 141
rect -311 107 -223 141
rect -133 107 -45 141
rect 45 107 133 141
rect 223 107 311 141
rect 401 107 489 141
rect 579 107 667 141
rect 757 107 845 141
<< locali >>
rect -1041 245 -945 279
rect 945 245 1041 279
rect -1041 183 -1007 245
rect 1007 183 1041 245
rect -861 107 -845 141
rect -757 107 -741 141
rect -683 107 -667 141
rect -579 107 -563 141
rect -505 107 -489 141
rect -401 107 -385 141
rect -327 107 -311 141
rect -223 107 -207 141
rect -149 107 -133 141
rect -45 107 -29 141
rect 29 107 45 141
rect 133 107 149 141
rect 207 107 223 141
rect 311 107 327 141
rect 385 107 401 141
rect 489 107 505 141
rect 563 107 579 141
rect 667 107 683 141
rect 741 107 757 141
rect 845 107 861 141
rect -907 57 -873 73
rect -907 -135 -873 -119
rect -729 57 -695 73
rect -729 -135 -695 -119
rect -551 57 -517 73
rect -551 -135 -517 -119
rect -373 57 -339 73
rect -373 -135 -339 -119
rect -195 57 -161 73
rect -195 -135 -161 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 161 57 195 73
rect 161 -135 195 -119
rect 339 57 373 73
rect 339 -135 373 -119
rect 517 57 551 73
rect 517 -135 551 -119
rect 695 57 729 73
rect 695 -135 729 -119
rect 873 57 907 73
rect 873 -135 907 -119
rect -1041 -245 -1007 -183
rect 1007 -245 1041 -183
rect -1041 -279 -945 -245
rect 945 -279 1041 -245
<< viali >>
rect -845 107 -757 141
rect -667 107 -579 141
rect -489 107 -401 141
rect -311 107 -223 141
rect -133 107 -45 141
rect 45 107 133 141
rect 223 107 311 141
rect 401 107 489 141
rect 579 107 667 141
rect 757 107 845 141
rect -907 -119 -873 57
rect -729 -119 -695 57
rect -551 -119 -517 57
rect -373 -119 -339 57
rect -195 -119 -161 57
rect -17 -119 17 57
rect 161 -119 195 57
rect 339 -119 373 57
rect 517 -119 551 57
rect 695 -119 729 57
rect 873 -119 907 57
<< metal1 >>
rect -857 141 -745 147
rect -857 107 -845 141
rect -757 107 -745 141
rect -857 101 -745 107
rect -679 141 -567 147
rect -679 107 -667 141
rect -579 107 -567 141
rect -679 101 -567 107
rect -501 141 -389 147
rect -501 107 -489 141
rect -401 107 -389 141
rect -501 101 -389 107
rect -323 141 -211 147
rect -323 107 -311 141
rect -223 107 -211 141
rect -323 101 -211 107
rect -145 141 -33 147
rect -145 107 -133 141
rect -45 107 -33 141
rect -145 101 -33 107
rect 33 141 145 147
rect 33 107 45 141
rect 133 107 145 141
rect 33 101 145 107
rect 211 141 323 147
rect 211 107 223 141
rect 311 107 323 141
rect 211 101 323 107
rect 389 141 501 147
rect 389 107 401 141
rect 489 107 501 141
rect 389 101 501 107
rect 567 141 679 147
rect 567 107 579 141
rect 667 107 679 141
rect 567 101 679 107
rect 745 141 857 147
rect 745 107 757 141
rect 845 107 857 141
rect 745 101 857 107
rect -913 57 -867 69
rect -913 -119 -907 57
rect -873 -119 -867 57
rect -913 -131 -867 -119
rect -735 57 -689 69
rect -735 -119 -729 57
rect -695 -119 -689 57
rect -735 -131 -689 -119
rect -557 57 -511 69
rect -557 -119 -551 57
rect -517 -119 -511 57
rect -557 -131 -511 -119
rect -379 57 -333 69
rect -379 -119 -373 57
rect -339 -119 -333 57
rect -379 -131 -333 -119
rect -201 57 -155 69
rect -201 -119 -195 57
rect -161 -119 -155 57
rect -201 -131 -155 -119
rect -23 57 23 69
rect -23 -119 -17 57
rect 17 -119 23 57
rect -23 -131 23 -119
rect 155 57 201 69
rect 155 -119 161 57
rect 195 -119 201 57
rect 155 -131 201 -119
rect 333 57 379 69
rect 333 -119 339 57
rect 373 -119 379 57
rect 333 -131 379 -119
rect 511 57 557 69
rect 511 -119 517 57
rect 551 -119 557 57
rect 511 -131 557 -119
rect 689 57 735 69
rect 689 -119 695 57
rect 729 -119 735 57
rect 689 -131 735 -119
rect 867 57 913 69
rect 867 -119 873 57
rect 907 -119 913 57
rect 867 -131 913 -119
<< properties >>
string FIXED_BBOX -1024 -262 1024 262
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.6 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
