magic
tech sky130A
magscale 1 2
timestamp 1712503184
<< error_s >>
rect -3924 4606 -3850 4615
rect -3924 4550 -3915 4606
rect -3924 4541 -3850 4550
rect -4407 4358 -4333 4367
rect -3924 4358 -3850 4367
rect -4407 4302 -4398 4358
rect -3924 4302 -3915 4358
rect -4407 4293 -4333 4302
rect -3924 4293 -3850 4302
rect 10492 -905 10618 -889
rect 11030 -1236 11083 -1086
rect 11191 -1401 11248 -1248
rect 11030 -1728 11083 -1578
rect 11030 -1938 11083 -1788
rect 11191 -1978 11248 -1413
rect 11030 -2143 11083 -2072
<< dnwell >>
rect -28958 10652 -6352 11020
rect -28958 499 -6351 10652
rect -28958 -5451 -10341 499
rect -28958 -16530 12219 -5451
<< nwell >>
rect -29038 10814 -6271 11100
rect -29038 -16324 -28752 10814
rect -6558 705 -6271 10814
rect -4967 707 -2959 761
rect -10547 419 -6271 705
rect -10547 -5371 -10261 419
rect -10547 -5657 12299 -5371
rect 12013 -16324 12299 -5657
rect -29038 -16610 12299 -16324
<< pwell >>
rect -4959 38 -2960 146
<< psubdiff >>
rect -4929 69 -4851 108
rect -3092 69 -2997 108
<< nsubdiff >>
rect -29001 11043 -6309 11063
rect -29001 11009 -28921 11043
rect -6415 11009 -6309 11043
rect -29001 10989 -6309 11009
rect -29001 10983 -28927 10989
rect -29001 -16493 -28981 10983
rect -28947 -16493 -28927 10983
rect -6383 10957 -6309 10989
rect -6383 536 -6363 10957
rect -6329 536 -6309 10957
rect -4929 686 -4870 725
rect -3070 686 -2997 725
rect -6383 530 -6309 536
rect -10372 510 -6309 530
rect -10372 476 -10292 510
rect -6389 476 -6309 510
rect -10372 456 -6309 476
rect -10372 449 -10298 456
rect -10372 -5328 -10352 449
rect -10318 -5328 -10298 449
rect -10372 -5408 -10298 -5328
rect -10372 -5428 12262 -5408
rect -10372 -5462 -10214 -5428
rect 12182 -5462 12262 -5428
rect -10372 -5482 12262 -5462
rect -29001 -16499 -28927 -16493
rect 12188 -5488 12262 -5482
rect 12188 -16493 12208 -5488
rect 12242 -16493 12262 -5488
rect 12188 -16499 12262 -16493
rect -29001 -16519 12262 -16499
rect -29001 -16553 -28921 -16519
rect 12182 -16553 12262 -16519
rect -29001 -16573 12262 -16553
<< psubdiffcont >>
rect -4851 69 -3092 108
<< nsubdiffcont >>
rect -28921 11009 -6415 11043
rect -28981 -16493 -28947 10983
rect -6363 536 -6329 10957
rect -4870 686 -3070 725
rect -10292 476 -6389 510
rect -10352 -5328 -10318 449
rect -10214 -5462 12182 -5428
rect 12208 -16493 12242 -5488
rect -28921 -16553 12182 -16519
<< locali >>
rect -28981 11009 -28921 11043
rect -6415 11009 -6329 11043
rect -28981 10983 -28947 11009
rect -6363 10957 -6329 11009
rect -15150 6793 -15086 6808
rect -15150 6695 -15135 6793
rect -15101 6695 -15086 6793
rect -15150 6680 -15086 6695
rect -4128 4664 -4000 4679
rect -4128 4566 -4113 4664
rect -4015 4566 -4000 4664
rect -3784 4664 -3720 4679
rect -4128 4551 -4000 4566
rect -3919 4595 -3855 4610
rect -3919 4561 -3904 4595
rect -3870 4561 -3855 4595
rect -3919 4546 -3855 4561
rect -3784 4566 -3769 4664
rect -3735 4566 -3720 4664
rect -3784 4551 -3720 4566
rect -3048 4548 -2990 4560
rect -3048 4514 -3036 4548
rect -3002 4514 -2990 4548
rect -3048 4502 -2990 4514
rect -3204 4406 -3076 4421
rect -3204 4308 -3189 4406
rect -3091 4308 -3076 4406
rect -2936 4406 -2872 4421
rect -3204 4293 -3076 4308
rect -3035 4342 -2971 4357
rect -3035 4308 -3020 4342
rect -2986 4308 -2971 4342
rect -3035 4293 -2971 4308
rect -2936 4308 -2921 4406
rect -2887 4308 -2872 4406
rect -2936 4293 -2872 4308
rect -3090 4038 -2962 4053
rect -3090 4004 -3075 4038
rect -2977 4004 -2962 4038
rect -3090 3989 -2962 4004
rect -4929 686 -4870 725
rect -3070 686 -2997 725
rect -6363 510 -6329 536
rect -10352 476 -10292 510
rect -6389 476 -6329 510
rect -10352 449 -10318 476
rect -4495 340 -4452 388
rect -3167 234 -3123 258
rect -4929 69 -4851 108
rect -3092 69 -2997 108
rect -6515 -1210 -6451 -1195
rect -6515 -1308 -6500 -1210
rect -6466 -1308 -6451 -1210
rect -6515 -1323 -6451 -1308
rect -4403 -1210 -4339 -1195
rect -4403 -1308 -4388 -1210
rect -4354 -1308 -4339 -1210
rect -4403 -1323 -4339 -1308
rect -2291 -1210 -2227 -1195
rect -2291 -1308 -2276 -1210
rect -2242 -1308 -2227 -1210
rect -2291 -1323 -2227 -1308
rect -179 -1210 -115 -1195
rect -179 -1308 -164 -1210
rect -130 -1308 -115 -1210
rect -179 -1323 -115 -1308
rect 1933 -1210 1997 -1195
rect 1933 -1308 1948 -1210
rect 1982 -1308 1997 -1210
rect 1933 -1323 1997 -1308
rect 4045 -1210 4109 -1195
rect 4045 -1308 4060 -1210
rect 4094 -1308 4109 -1210
rect 4045 -1323 4109 -1308
rect 6157 -1210 6221 -1195
rect 6157 -1308 6172 -1210
rect 6206 -1308 6221 -1210
rect 6157 -1323 6221 -1308
rect 8269 -1210 8333 -1195
rect 8269 -1308 8284 -1210
rect 8318 -1308 8333 -1210
rect 8269 -1323 8333 -1308
rect 10381 -1210 10445 -1195
rect 10381 -1308 10396 -1210
rect 10430 -1308 10445 -1210
rect 10381 -1323 10445 -1308
rect 11174 -1843 11250 -1831
rect 11174 -1895 11186 -1843
rect 11238 -1895 11250 -1843
rect 11174 -1907 11250 -1895
rect -8047 -1942 -7983 -1927
rect -8047 -2040 -8032 -1942
rect -7998 -2040 -7983 -1942
rect -8047 -2055 -7983 -2040
rect -5935 -1942 -5871 -1927
rect -5935 -2040 -5920 -1942
rect -5886 -2040 -5871 -1942
rect -5935 -2055 -5871 -2040
rect -3823 -1942 -3759 -1927
rect -3823 -2040 -3808 -1942
rect -3774 -2040 -3759 -1942
rect -3823 -2055 -3759 -2040
rect -1711 -1942 -1647 -1927
rect -1711 -2040 -1696 -1942
rect -1662 -2040 -1647 -1942
rect -1711 -2055 -1647 -2040
rect 401 -1942 465 -1927
rect 401 -2040 416 -1942
rect 450 -2040 465 -1942
rect 401 -2055 465 -2040
rect 2513 -1942 2577 -1927
rect 2513 -2040 2528 -1942
rect 2562 -2040 2577 -1942
rect 2513 -2055 2577 -2040
rect 4625 -1942 4689 -1927
rect 4625 -2040 4640 -1942
rect 4674 -2040 4689 -1942
rect 4625 -2055 4689 -2040
rect 6737 -1942 6801 -1927
rect 6737 -2040 6752 -1942
rect 6786 -2040 6801 -1942
rect 6737 -2055 6801 -2040
rect 8849 -1942 8913 -1927
rect 8849 -2040 8864 -1942
rect 8898 -2040 8913 -1942
rect 8849 -2055 8913 -2040
rect -6515 -2944 -6451 -2929
rect -6515 -3042 -6500 -2944
rect -6466 -3042 -6451 -2944
rect -6515 -3057 -6451 -3042
rect -4403 -2944 -4339 -2929
rect -4403 -3042 -4388 -2944
rect -4354 -3042 -4339 -2944
rect -4403 -3057 -4339 -3042
rect -2291 -2944 -2227 -2929
rect -2291 -3042 -2276 -2944
rect -2242 -3042 -2227 -2944
rect -2291 -3057 -2227 -3042
rect -179 -2944 -115 -2929
rect -179 -3042 -164 -2944
rect -130 -3042 -115 -2944
rect -179 -3057 -115 -3042
rect 1933 -2944 1997 -2929
rect 1933 -3042 1948 -2944
rect 1982 -3042 1997 -2944
rect 1933 -3057 1997 -3042
rect 4045 -2944 4109 -2929
rect 4045 -3042 4060 -2944
rect 4094 -3042 4109 -2944
rect 4045 -3057 4109 -3042
rect 6157 -2944 6221 -2929
rect 6157 -3042 6172 -2944
rect 6206 -3042 6221 -2944
rect 6157 -3057 6221 -3042
rect 8269 -2944 8333 -2929
rect 8269 -3042 8284 -2944
rect 8318 -3042 8333 -2944
rect 8269 -3057 8333 -3042
rect 10381 -2944 10445 -2929
rect 10381 -3042 10396 -2944
rect 10430 -3042 10445 -2944
rect 10381 -3057 10445 -3042
rect -8047 -3676 -7983 -3661
rect -8047 -3774 -8032 -3676
rect -7998 -3774 -7983 -3676
rect -8047 -3789 -7983 -3774
rect -5935 -3676 -5871 -3661
rect -5935 -3774 -5920 -3676
rect -5886 -3774 -5871 -3676
rect -5935 -3789 -5871 -3774
rect -3823 -3676 -3759 -3661
rect -3823 -3774 -3808 -3676
rect -3774 -3774 -3759 -3676
rect -3823 -3789 -3759 -3774
rect -1711 -3676 -1647 -3661
rect -1711 -3774 -1696 -3676
rect -1662 -3774 -1647 -3676
rect -1711 -3789 -1647 -3774
rect 401 -3676 465 -3661
rect 401 -3774 416 -3676
rect 450 -3774 465 -3676
rect 401 -3789 465 -3774
rect 2513 -3676 2577 -3661
rect 2513 -3774 2528 -3676
rect 2562 -3774 2577 -3676
rect 2513 -3789 2577 -3774
rect 4625 -3676 4689 -3661
rect 4625 -3774 4640 -3676
rect 4674 -3774 4689 -3676
rect 4625 -3789 4689 -3774
rect 6737 -3676 6801 -3661
rect 6737 -3774 6752 -3676
rect 6786 -3774 6801 -3676
rect 6737 -3789 6801 -3774
rect 8849 -3676 8913 -3661
rect 8849 -3774 8864 -3676
rect 8898 -3774 8913 -3676
rect 8849 -3789 8913 -3774
rect -10352 -5428 -10318 -5328
rect -10352 -5462 -10214 -5428
rect 12182 -5462 12242 -5428
rect 12208 -5488 12242 -5462
rect -28981 -16519 -28947 -16493
rect 12208 -16519 12242 -16493
rect -28981 -16553 -28921 -16519
rect 12182 -16553 12242 -16519
<< viali >>
rect -29003 10119 -28981 10255
rect -28981 10119 -28947 10255
rect -28947 10119 -28867 10255
rect -15135 6695 -15101 6793
rect -4113 4566 -4015 4664
rect -3904 4561 -3870 4595
rect -3769 4566 -3735 4664
rect -3036 4514 -3002 4548
rect -3189 4308 -3091 4406
rect -3020 4308 -2986 4342
rect -2921 4308 -2887 4406
rect -3075 4004 -2977 4038
rect -4888 346 -4644 380
rect -3167 258 -3123 495
rect -6500 -1308 -6466 -1210
rect -4388 -1308 -4354 -1210
rect -2276 -1308 -2242 -1210
rect -164 -1308 -130 -1210
rect 1948 -1308 1982 -1210
rect 4060 -1308 4094 -1210
rect 6172 -1308 6206 -1210
rect 8284 -1308 8318 -1210
rect 10396 -1308 10430 -1210
rect 10642 -1378 10690 -1330
rect 11186 -1895 11238 -1843
rect -8032 -2040 -7998 -1942
rect -5920 -2040 -5886 -1942
rect -3808 -2040 -3774 -1942
rect -1696 -2040 -1662 -1942
rect 416 -2040 450 -1942
rect 2528 -2040 2562 -1942
rect 4640 -2040 4674 -1942
rect 6752 -2040 6786 -1942
rect 8864 -2040 8898 -1942
rect -6500 -3042 -6466 -2944
rect -4388 -3042 -4354 -2944
rect -2276 -3042 -2242 -2944
rect -164 -3042 -130 -2944
rect 1948 -3042 1982 -2944
rect 4060 -3042 4094 -2944
rect 6172 -3042 6206 -2944
rect 8284 -3042 8318 -2944
rect 10396 -3042 10430 -2944
rect -8032 -3774 -7998 -3676
rect -5920 -3774 -5886 -3676
rect -3808 -3774 -3774 -3676
rect -1696 -3774 -1662 -3676
rect 416 -3774 450 -3676
rect 2528 -3774 2562 -3676
rect 4640 -3774 4674 -3676
rect 6752 -3774 6786 -3676
rect 8864 -3774 8898 -3676
rect -29009 -11096 -28981 -10858
rect -28981 -11096 -28947 -10858
rect -28947 -11096 -28771 -10858
<< metal1 >>
rect -29015 10261 -28855 10267
rect -29015 10113 -29009 10261
rect -28861 10113 -28855 10261
rect -29015 10107 -28855 10113
rect -14727 9400 -14611 9821
rect -13971 9400 -13855 9821
rect -13215 9400 -13099 9821
rect -12459 9400 -12343 9821
rect -11703 9400 -11587 9821
rect -10947 9400 -10831 9821
rect -10191 9400 -10075 9821
rect -9435 9400 -9319 9821
rect -8679 9400 -8563 9821
rect -7923 9400 -7807 9821
rect -15155 6807 -15081 6818
rect -15155 6681 -15144 6807
rect -15092 6681 -15081 6807
rect -15155 6670 -15081 6681
rect -4138 4678 -3990 4689
rect -4138 4552 -4127 4678
rect -4001 4552 -3990 4678
rect -3789 4678 -3715 4689
rect -4138 4541 -3990 4552
rect -3924 4604 -3850 4615
rect -3924 4552 -3913 4604
rect -3861 4552 -3850 4604
rect -3924 4541 -3850 4552
rect -3789 4552 -3778 4678
rect -3726 4552 -3715 4678
rect -3789 4541 -3715 4552
rect -3048 4548 -2990 4560
rect -3048 4514 -3036 4548
rect -3002 4514 -2990 4548
rect -3048 4502 -2990 4514
rect -4138 4430 -3990 4441
rect -4138 4304 -4127 4430
rect -4001 4304 -3990 4430
rect -3789 4430 -3715 4441
rect -4138 4293 -3990 4304
rect -3924 4356 -3850 4367
rect -3924 4304 -3913 4356
rect -3861 4304 -3850 4356
rect -3924 4293 -3850 4304
rect -3789 4304 -3778 4430
rect -3726 4304 -3715 4430
rect -3789 4293 -3715 4304
rect -3632 4415 -3504 4421
rect -3632 4299 -3626 4415
rect -3510 4299 -3504 4415
rect -3364 4415 -3300 4421
rect -3632 4293 -3504 4299
rect -3463 4351 -3399 4357
rect -3463 4299 -3457 4351
rect -3405 4299 -3399 4351
rect -3463 4293 -3399 4299
rect -3364 4299 -3358 4415
rect -3306 4299 -3300 4415
rect -3364 4293 -3300 4299
rect -3204 4415 -3076 4421
rect -3204 4299 -3198 4415
rect -3082 4299 -3076 4415
rect -2936 4415 -2872 4421
rect -3204 4293 -3076 4299
rect -3035 4351 -2971 4357
rect -3035 4299 -3029 4351
rect -2977 4299 -2971 4351
rect -3035 4293 -2971 4299
rect -2936 4299 -2930 4415
rect -2878 4299 -2872 4415
rect -2936 4293 -2872 4299
rect -3344 4121 -3216 4127
rect -3344 4069 -3338 4121
rect -3222 4069 -3216 4121
rect -3344 4063 -3216 4069
rect -3090 4047 -2962 4053
rect -3780 4032 -3632 4043
rect -3780 3980 -3769 4032
rect -3643 3980 -3632 4032
rect -3090 3995 -3084 4047
rect -2968 3995 -2962 4047
rect -3090 3989 -2962 3995
rect -3780 3969 -3632 3980
rect -14892 2029 -14886 2093
rect -14822 2029 -14816 2093
rect -14349 2001 -14233 2422
rect -13593 2001 -13477 2422
rect -12837 2001 -12721 2422
rect -12081 2001 -11965 2422
rect -11325 2001 -11209 2422
rect -10569 2001 -10453 2422
rect -9813 2001 -9697 2422
rect -9057 2001 -8941 2422
rect -8301 2001 -8185 2422
rect -7731 2013 -7725 2107
rect -7621 2013 -7615 2107
rect -5486 2042 -5027 2048
rect -5486 1883 -5478 2042
rect -5364 1883 -5027 2042
rect -5486 1876 -5027 1883
rect -5286 1397 -4999 1402
rect -5286 1240 -5277 1397
rect -5167 1240 -4999 1397
rect -5286 1233 -4999 1240
rect -5486 706 -4929 717
rect -5486 630 -5477 706
rect -5370 630 -4929 706
rect -5486 621 -4929 630
rect -3173 496 -3117 508
rect -4903 380 -4696 395
rect -4903 346 -4888 380
rect -4903 335 -4696 346
rect -4636 335 -4630 395
rect -3173 228 -3117 241
rect -5286 167 -4929 173
rect -5286 83 -5278 167
rect -5166 83 -4929 167
rect -5286 77 -4929 83
rect -9258 -593 -9252 -465
rect -9124 -593 -5486 -465
rect -5358 -593 -5352 -465
rect -8852 -718 -6055 -712
rect -8852 -854 -8846 -718
rect -8730 -724 -6055 -718
rect -5918 -724 11768 -712
rect -8730 -732 11768 -724
rect -8730 -854 -5286 -732
rect -8852 -860 -5286 -854
rect -5158 -860 11768 -732
rect -6515 -1201 -6451 -1195
rect -6515 -1317 -6509 -1201
rect -6457 -1317 -6451 -1201
rect -6515 -1323 -6451 -1317
rect -4403 -1201 -4339 -1195
rect -4403 -1317 -4397 -1201
rect -4345 -1317 -4339 -1201
rect -4403 -1323 -4339 -1317
rect -2291 -1201 -2227 -1195
rect -2291 -1317 -2285 -1201
rect -2233 -1317 -2227 -1201
rect -2291 -1323 -2227 -1317
rect -179 -1201 -115 -1195
rect -179 -1317 -173 -1201
rect -121 -1317 -115 -1201
rect -179 -1323 -115 -1317
rect 1933 -1201 1997 -1195
rect 1933 -1317 1939 -1201
rect 1991 -1317 1997 -1201
rect 1933 -1323 1997 -1317
rect 4045 -1201 4109 -1195
rect 4045 -1317 4051 -1201
rect 4103 -1317 4109 -1201
rect 4045 -1323 4109 -1317
rect 6157 -1201 6221 -1195
rect 6157 -1317 6163 -1201
rect 6215 -1317 6221 -1201
rect 6157 -1323 6221 -1317
rect 8269 -1201 8333 -1195
rect 8269 -1317 8275 -1201
rect 8327 -1317 8333 -1201
rect 8269 -1323 8333 -1317
rect 10381 -1201 10445 -1195
rect 10381 -1317 10387 -1201
rect 10439 -1317 10445 -1201
rect 10381 -1323 10445 -1317
rect 10630 -1384 10636 -1324
rect 10696 -1384 10702 -1324
rect -9052 -1430 11768 -1424
rect -9052 -1668 -9046 -1430
rect -8930 -1668 11768 -1430
rect -9052 -1674 11768 -1668
rect -9252 -1704 12099 -1702
rect -9252 -1756 -9246 -1704
rect -9130 -1756 12099 -1704
rect -9252 -1759 12099 -1756
rect 11174 -1837 11250 -1831
rect 11174 -1901 11180 -1837
rect 11244 -1901 11250 -1837
rect 11174 -1907 11250 -1901
rect -8047 -1933 -7983 -1927
rect -8047 -2049 -8041 -1933
rect -7989 -2049 -7983 -1933
rect -8047 -2055 -7983 -2049
rect -5935 -1933 -5871 -1927
rect -5935 -2049 -5929 -1933
rect -5877 -2049 -5871 -1933
rect -5935 -2055 -5871 -2049
rect -3823 -1933 -3759 -1927
rect -3823 -2049 -3817 -1933
rect -3765 -2049 -3759 -1933
rect -3823 -2055 -3759 -2049
rect -1711 -1933 -1647 -1927
rect -1711 -2049 -1705 -1933
rect -1653 -2049 -1647 -1933
rect -1711 -2055 -1647 -2049
rect 401 -1933 465 -1927
rect 401 -2049 407 -1933
rect 459 -2049 465 -1933
rect 401 -2055 465 -2049
rect 2513 -1933 2577 -1927
rect 2513 -2049 2519 -1933
rect 2571 -2049 2577 -1933
rect 2513 -2055 2577 -2049
rect 4625 -1933 4689 -1927
rect 4625 -2049 4631 -1933
rect 4683 -2049 4689 -1933
rect 4625 -2055 4689 -2049
rect 6737 -1933 6801 -1927
rect 6737 -2049 6743 -1933
rect 6795 -2049 6801 -1933
rect 6737 -2055 6801 -2049
rect 8849 -1933 8913 -1927
rect 8849 -2049 8855 -1933
rect 8907 -2049 8913 -1933
rect 8849 -2055 8913 -2049
rect -8852 -2244 11768 -2238
rect -8852 -2588 -8846 -2244
rect -8730 -2588 11768 -2244
rect -8852 -2594 11768 -2588
rect -6515 -2935 -6451 -2929
rect -6515 -3051 -6509 -2935
rect -6457 -3051 -6451 -2935
rect -6515 -3057 -6451 -3051
rect -4403 -2935 -4339 -2929
rect -4403 -3051 -4397 -2935
rect -4345 -3051 -4339 -2935
rect -4403 -3057 -4339 -3051
rect -2291 -2935 -2227 -2929
rect -2291 -3051 -2285 -2935
rect -2233 -3051 -2227 -2935
rect -2291 -3057 -2227 -3051
rect -179 -2935 -115 -2929
rect -179 -3051 -173 -2935
rect -121 -3051 -115 -2935
rect -179 -3057 -115 -3051
rect 1933 -2935 1997 -2929
rect 1933 -3051 1939 -2935
rect 1991 -3051 1997 -2935
rect 1933 -3057 1997 -3051
rect 4045 -2935 4109 -2929
rect 4045 -3051 4051 -2935
rect 4103 -3051 4109 -2935
rect 4045 -3057 4109 -3051
rect 6157 -2935 6221 -2929
rect 6157 -3051 6163 -2935
rect 6215 -3051 6221 -2935
rect 6157 -3057 6221 -3051
rect 8269 -2935 8333 -2929
rect 8269 -3051 8275 -2935
rect 8327 -3051 8333 -2935
rect 8269 -3057 8333 -3051
rect 10381 -2935 10445 -2929
rect 10381 -3051 10387 -2935
rect 10439 -3051 10445 -2935
rect 10381 -3057 10445 -3051
rect -9052 -3164 10468 -3158
rect -9052 -3402 -9046 -3164
rect -8930 -3402 10468 -3164
rect -9052 -3408 10468 -3402
rect -9252 -3438 10471 -3436
rect -9252 -3490 -9246 -3438
rect -9130 -3490 10471 -3438
rect -9252 -3493 10471 -3490
rect -8047 -3667 -7983 -3661
rect -8047 -3783 -8041 -3667
rect -7989 -3783 -7983 -3667
rect -8047 -3789 -7983 -3783
rect -5935 -3667 -5871 -3661
rect -5935 -3783 -5929 -3667
rect -5877 -3783 -5871 -3667
rect -5935 -3789 -5871 -3783
rect -3823 -3667 -3759 -3661
rect -3823 -3783 -3817 -3667
rect -3765 -3783 -3759 -3667
rect -3823 -3789 -3759 -3783
rect -1711 -3667 -1647 -3661
rect -1711 -3783 -1705 -3667
rect -1653 -3783 -1647 -3667
rect -1711 -3789 -1647 -3783
rect 401 -3667 465 -3661
rect 401 -3783 407 -3667
rect 459 -3783 465 -3667
rect 401 -3789 465 -3783
rect 2513 -3667 2577 -3661
rect 2513 -3783 2519 -3667
rect 2571 -3783 2577 -3667
rect 2513 -3789 2577 -3783
rect 4625 -3667 4689 -3661
rect 4625 -3783 4631 -3667
rect 4683 -3783 4689 -3667
rect 4625 -3789 4689 -3783
rect 6737 -3667 6801 -3661
rect 6737 -3783 6743 -3667
rect 6795 -3783 6801 -3667
rect 6737 -3789 6801 -3783
rect 8849 -3667 8913 -3661
rect 8849 -3783 8855 -3667
rect 8907 -3783 8913 -3667
rect 8849 -3789 8913 -3783
rect -8852 -3978 10468 -3972
rect -8852 -4082 -8846 -3978
rect -9252 -4114 -8846 -4082
rect -8730 -4114 10468 -3978
rect -9252 -4282 10468 -4114
rect -9252 -4344 10468 -4338
rect -9252 -4532 -9246 -4344
rect -9130 -4532 10468 -4344
rect -9252 -4538 10468 -4532
rect -9252 -4600 10468 -4594
rect -9252 -4788 -9046 -4600
rect -8930 -4788 10468 -4600
rect -9252 -4794 10468 -4788
rect -4837 -6994 -4637 -4794
rect -27806 -10519 -27406 -10513
rect -27806 -10796 -27800 -10519
rect -27412 -10796 -27406 -10519
rect -27806 -10802 -27406 -10796
rect -19274 -10802 -10164 -10552
rect -10355 -10824 -10164 -10802
rect -10355 -10830 -4887 -10824
rect -29021 -10858 -27459 -10852
rect -29021 -11096 -29009 -10858
rect -28771 -11096 -28256 -10858
rect -27868 -11096 -27459 -10858
rect -29021 -11102 -27459 -11096
rect -19020 -11080 -10420 -10854
rect -10355 -11018 -5076 -10830
rect -4893 -11018 -4887 -10830
rect -10355 -11024 -4887 -11018
rect -19020 -11104 -4637 -11080
rect -10614 -11280 -4637 -11104
<< via1 >>
rect -29009 10255 -28861 10261
rect -29009 10119 -29003 10255
rect -29003 10119 -28867 10255
rect -28867 10119 -28861 10255
rect -29009 10113 -28861 10119
rect -15144 6793 -15092 6807
rect -15144 6695 -15135 6793
rect -15135 6695 -15101 6793
rect -15101 6695 -15092 6793
rect -15144 6681 -15092 6695
rect -4127 4664 -4001 4678
rect -4127 4566 -4113 4664
rect -4113 4566 -4015 4664
rect -4015 4566 -4001 4664
rect -4127 4552 -4001 4566
rect -3913 4595 -3861 4604
rect -3913 4561 -3904 4595
rect -3904 4561 -3870 4595
rect -3870 4561 -3861 4595
rect -3913 4552 -3861 4561
rect -3778 4664 -3726 4678
rect -3778 4566 -3769 4664
rect -3769 4566 -3735 4664
rect -3735 4566 -3726 4664
rect -3778 4552 -3726 4566
rect -4127 4304 -4001 4430
rect -3913 4304 -3861 4356
rect -3778 4304 -3726 4430
rect -3626 4299 -3510 4415
rect -3457 4299 -3405 4351
rect -3358 4299 -3306 4415
rect -3198 4406 -3082 4415
rect -3198 4308 -3189 4406
rect -3189 4308 -3091 4406
rect -3091 4308 -3082 4406
rect -3198 4299 -3082 4308
rect -3029 4342 -2977 4351
rect -3029 4308 -3020 4342
rect -3020 4308 -2986 4342
rect -2986 4308 -2977 4342
rect -3029 4299 -2977 4308
rect -2930 4406 -2878 4415
rect -2930 4308 -2921 4406
rect -2921 4308 -2887 4406
rect -2887 4308 -2878 4406
rect -2930 4299 -2878 4308
rect -3338 4069 -3222 4121
rect -3769 3980 -3643 4032
rect -3084 4038 -2968 4047
rect -3084 4004 -3075 4038
rect -3075 4004 -2977 4038
rect -2977 4004 -2968 4038
rect -3084 3995 -2968 4004
rect -14886 2029 -14822 2093
rect -7725 2013 -7621 2107
rect -5478 1883 -5364 2042
rect -5277 1240 -5167 1397
rect -5477 630 -5370 706
rect -3173 495 -3117 496
rect -4696 380 -4636 395
rect -4696 346 -4644 380
rect -4644 346 -4636 380
rect -4696 335 -4636 346
rect -3173 258 -3167 495
rect -3167 258 -3123 495
rect -3123 258 -3117 495
rect -3173 241 -3117 258
rect -5278 83 -5166 167
rect -9252 -593 -9124 -465
rect -5486 -593 -5358 -465
rect -8846 -854 -8730 -718
rect -5286 -860 -5158 -732
rect -6509 -1210 -6457 -1201
rect -6509 -1308 -6500 -1210
rect -6500 -1308 -6466 -1210
rect -6466 -1308 -6457 -1210
rect -6509 -1317 -6457 -1308
rect -4397 -1210 -4345 -1201
rect -4397 -1308 -4388 -1210
rect -4388 -1308 -4354 -1210
rect -4354 -1308 -4345 -1210
rect -4397 -1317 -4345 -1308
rect -2285 -1210 -2233 -1201
rect -2285 -1308 -2276 -1210
rect -2276 -1308 -2242 -1210
rect -2242 -1308 -2233 -1210
rect -2285 -1317 -2233 -1308
rect -173 -1210 -121 -1201
rect -173 -1308 -164 -1210
rect -164 -1308 -130 -1210
rect -130 -1308 -121 -1210
rect -173 -1317 -121 -1308
rect 1939 -1210 1991 -1201
rect 1939 -1308 1948 -1210
rect 1948 -1308 1982 -1210
rect 1982 -1308 1991 -1210
rect 1939 -1317 1991 -1308
rect 4051 -1210 4103 -1201
rect 4051 -1308 4060 -1210
rect 4060 -1308 4094 -1210
rect 4094 -1308 4103 -1210
rect 4051 -1317 4103 -1308
rect 6163 -1210 6215 -1201
rect 6163 -1308 6172 -1210
rect 6172 -1308 6206 -1210
rect 6206 -1308 6215 -1210
rect 6163 -1317 6215 -1308
rect 8275 -1210 8327 -1201
rect 8275 -1308 8284 -1210
rect 8284 -1308 8318 -1210
rect 8318 -1308 8327 -1210
rect 8275 -1317 8327 -1308
rect 10387 -1210 10439 -1201
rect 10387 -1308 10396 -1210
rect 10396 -1308 10430 -1210
rect 10430 -1308 10439 -1210
rect 10387 -1317 10439 -1308
rect 10636 -1330 10696 -1324
rect 10636 -1378 10642 -1330
rect 10642 -1378 10690 -1330
rect 10690 -1378 10696 -1330
rect 10636 -1384 10696 -1378
rect -9046 -1668 -8930 -1430
rect -9246 -1756 -9130 -1704
rect 11180 -1843 11244 -1837
rect 11180 -1895 11186 -1843
rect 11186 -1895 11238 -1843
rect 11238 -1895 11244 -1843
rect 11180 -1901 11244 -1895
rect -8041 -1942 -7989 -1933
rect -8041 -2040 -8032 -1942
rect -8032 -2040 -7998 -1942
rect -7998 -2040 -7989 -1942
rect -8041 -2049 -7989 -2040
rect -5929 -1942 -5877 -1933
rect -5929 -2040 -5920 -1942
rect -5920 -2040 -5886 -1942
rect -5886 -2040 -5877 -1942
rect -5929 -2049 -5877 -2040
rect -3817 -1942 -3765 -1933
rect -3817 -2040 -3808 -1942
rect -3808 -2040 -3774 -1942
rect -3774 -2040 -3765 -1942
rect -3817 -2049 -3765 -2040
rect -1705 -1942 -1653 -1933
rect -1705 -2040 -1696 -1942
rect -1696 -2040 -1662 -1942
rect -1662 -2040 -1653 -1942
rect -1705 -2049 -1653 -2040
rect 407 -1942 459 -1933
rect 407 -2040 416 -1942
rect 416 -2040 450 -1942
rect 450 -2040 459 -1942
rect 407 -2049 459 -2040
rect 2519 -1942 2571 -1933
rect 2519 -2040 2528 -1942
rect 2528 -2040 2562 -1942
rect 2562 -2040 2571 -1942
rect 2519 -2049 2571 -2040
rect 4631 -1942 4683 -1933
rect 4631 -2040 4640 -1942
rect 4640 -2040 4674 -1942
rect 4674 -2040 4683 -1942
rect 4631 -2049 4683 -2040
rect 6743 -1942 6795 -1933
rect 6743 -2040 6752 -1942
rect 6752 -2040 6786 -1942
rect 6786 -2040 6795 -1942
rect 6743 -2049 6795 -2040
rect 8855 -1942 8907 -1933
rect 8855 -2040 8864 -1942
rect 8864 -2040 8898 -1942
rect 8898 -2040 8907 -1942
rect 8855 -2049 8907 -2040
rect -8846 -2588 -8730 -2244
rect -6509 -2944 -6457 -2935
rect -6509 -3042 -6500 -2944
rect -6500 -3042 -6466 -2944
rect -6466 -3042 -6457 -2944
rect -6509 -3051 -6457 -3042
rect -4397 -2944 -4345 -2935
rect -4397 -3042 -4388 -2944
rect -4388 -3042 -4354 -2944
rect -4354 -3042 -4345 -2944
rect -4397 -3051 -4345 -3042
rect -2285 -2944 -2233 -2935
rect -2285 -3042 -2276 -2944
rect -2276 -3042 -2242 -2944
rect -2242 -3042 -2233 -2944
rect -2285 -3051 -2233 -3042
rect -173 -2944 -121 -2935
rect -173 -3042 -164 -2944
rect -164 -3042 -130 -2944
rect -130 -3042 -121 -2944
rect -173 -3051 -121 -3042
rect 1939 -2944 1991 -2935
rect 1939 -3042 1948 -2944
rect 1948 -3042 1982 -2944
rect 1982 -3042 1991 -2944
rect 1939 -3051 1991 -3042
rect 4051 -2944 4103 -2935
rect 4051 -3042 4060 -2944
rect 4060 -3042 4094 -2944
rect 4094 -3042 4103 -2944
rect 4051 -3051 4103 -3042
rect 6163 -2944 6215 -2935
rect 6163 -3042 6172 -2944
rect 6172 -3042 6206 -2944
rect 6206 -3042 6215 -2944
rect 6163 -3051 6215 -3042
rect 8275 -2944 8327 -2935
rect 8275 -3042 8284 -2944
rect 8284 -3042 8318 -2944
rect 8318 -3042 8327 -2944
rect 8275 -3051 8327 -3042
rect 10387 -2944 10439 -2935
rect 10387 -3042 10396 -2944
rect 10396 -3042 10430 -2944
rect 10430 -3042 10439 -2944
rect 10387 -3051 10439 -3042
rect -9046 -3402 -8930 -3164
rect -9246 -3490 -9130 -3438
rect -8041 -3676 -7989 -3667
rect -8041 -3774 -8032 -3676
rect -8032 -3774 -7998 -3676
rect -7998 -3774 -7989 -3676
rect -8041 -3783 -7989 -3774
rect -5929 -3676 -5877 -3667
rect -5929 -3774 -5920 -3676
rect -5920 -3774 -5886 -3676
rect -5886 -3774 -5877 -3676
rect -5929 -3783 -5877 -3774
rect -3817 -3676 -3765 -3667
rect -3817 -3774 -3808 -3676
rect -3808 -3774 -3774 -3676
rect -3774 -3774 -3765 -3676
rect -3817 -3783 -3765 -3774
rect -1705 -3676 -1653 -3667
rect -1705 -3774 -1696 -3676
rect -1696 -3774 -1662 -3676
rect -1662 -3774 -1653 -3676
rect -1705 -3783 -1653 -3774
rect 407 -3676 459 -3667
rect 407 -3774 416 -3676
rect 416 -3774 450 -3676
rect 450 -3774 459 -3676
rect 407 -3783 459 -3774
rect 2519 -3676 2571 -3667
rect 2519 -3774 2528 -3676
rect 2528 -3774 2562 -3676
rect 2562 -3774 2571 -3676
rect 2519 -3783 2571 -3774
rect 4631 -3676 4683 -3667
rect 4631 -3774 4640 -3676
rect 4640 -3774 4674 -3676
rect 4674 -3774 4683 -3676
rect 4631 -3783 4683 -3774
rect 6743 -3676 6795 -3667
rect 6743 -3774 6752 -3676
rect 6752 -3774 6786 -3676
rect 6786 -3774 6795 -3676
rect 6743 -3783 6795 -3774
rect 8855 -3676 8907 -3667
rect 8855 -3774 8864 -3676
rect 8864 -3774 8898 -3676
rect 8898 -3774 8907 -3676
rect 8855 -3783 8907 -3774
rect -8846 -4114 -8730 -3978
rect -9246 -4532 -9130 -4344
rect -9046 -4788 -8930 -4600
rect -27800 -10796 -27412 -10519
rect -28256 -11096 -27868 -10858
rect -5076 -11018 -4893 -10830
rect -4575 -11018 -4387 -10830
<< metal2 >>
rect -29015 10261 -28855 10267
rect -29015 10113 -29009 10261
rect -28861 10113 -28855 10261
rect -29015 10107 -28855 10113
rect -28262 10255 -27862 10398
rect -28262 10119 -27929 10255
rect -27868 10119 -27862 10255
rect -29931 -1228 -29793 -1224
rect -29936 -1233 -29788 -1228
rect -29936 -1371 -29931 -1233
rect -29793 -1371 -29788 -1233
rect -29936 -1534 -29788 -1371
rect -28262 -10858 -27862 10119
rect -27806 6812 -27406 10398
rect -19249 7756 -19185 7760
rect -19254 7751 -19180 7756
rect -19254 7687 -19249 7751
rect -19185 7687 -19180 7751
rect -27035 7147 -26979 7156
rect -27035 7082 -26979 7091
rect -27806 6676 -27478 6812
rect -27412 6676 -27406 6812
rect -27806 2314 -27406 6676
rect -27806 2178 -27478 2314
rect -27412 2178 -27406 2314
rect -27806 -10519 -27406 2178
rect -19254 607 -19180 7687
rect -17661 7151 -17597 7160
rect -18588 5514 -18528 5523
rect -18588 -8044 -18528 5454
rect -18293 5314 -18229 5323
rect -18293 2438 -18229 5250
rect -18293 2374 -18177 2438
rect -18241 -2878 -18177 2374
rect -17661 -2678 -17597 7087
rect -17531 605 -17457 753
rect -16331 -763 -16275 7374
rect -15155 6809 -15081 6818
rect -15155 6679 -15146 6809
rect -15090 6679 -15081 6809
rect -15155 6670 -15081 6679
rect -4138 4680 -3990 4689
rect -4138 4550 -4129 4680
rect -3999 4550 -3990 4680
rect -3789 4680 -3715 4689
rect -4138 4541 -3990 4550
rect -3924 4606 -3850 4615
rect -3924 4550 -3915 4606
rect -3859 4550 -3850 4606
rect -3924 4541 -3850 4550
rect -3789 4550 -3780 4680
rect -3724 4550 -3715 4680
rect -3789 4541 -3715 4550
rect -4622 4432 -4474 4441
rect -4622 4302 -4613 4432
rect -4483 4302 -4474 4432
rect -4273 4432 -4199 4441
rect -4622 4293 -4474 4302
rect -4407 4358 -4333 4367
rect -4407 4302 -4398 4358
rect -4342 4302 -4333 4358
rect -4407 4293 -4333 4302
rect -4273 4302 -4264 4432
rect -4208 4302 -4199 4432
rect -4273 4293 -4199 4302
rect -4138 4432 -3990 4441
rect -4138 4302 -4129 4432
rect -3999 4302 -3990 4432
rect -3789 4432 -3715 4441
rect -4138 4293 -3990 4302
rect -3924 4358 -3850 4367
rect -3924 4302 -3915 4358
rect -3859 4302 -3850 4358
rect -3924 4293 -3850 4302
rect -3789 4302 -3780 4432
rect -3724 4302 -3715 4432
rect -3789 4293 -3715 4302
rect -3632 4415 -3504 4421
rect -3632 4299 -3626 4415
rect -3510 4299 -3504 4415
rect -3364 4415 -3300 4421
rect -3632 4293 -3504 4299
rect -3463 4351 -3399 4357
rect -3463 4299 -3457 4351
rect -3405 4299 -3399 4351
rect -3463 4293 -3399 4299
rect -3364 4299 -3358 4415
rect -3306 4299 -3300 4415
rect -3364 4293 -3300 4299
rect -3204 4415 -3076 4421
rect -3204 4299 -3198 4415
rect -3082 4299 -3076 4415
rect -2936 4415 -2872 4421
rect -3204 4293 -3076 4299
rect -3035 4351 -2971 4357
rect -3035 4299 -3029 4351
rect -2977 4299 -2971 4351
rect -3035 4293 -2971 4299
rect -2936 4299 -2930 4415
rect -2878 4299 -2872 4415
rect -2936 4293 -2872 4299
rect -3344 4121 -3216 4127
rect -4264 4078 -4116 4087
rect -4264 4022 -4255 4078
rect -4125 4022 -4116 4078
rect -3344 4069 -3338 4121
rect -3222 4069 -3216 4121
rect -3344 4063 -3216 4069
rect -3090 4047 -2962 4053
rect -4264 4013 -4116 4022
rect -3780 4034 -3632 4043
rect -3780 3978 -3771 4034
rect -3641 3978 -3632 4034
rect -3090 3995 -3084 4047
rect -2968 3995 -2962 4047
rect -3090 3989 -2962 3995
rect -3780 3969 -3632 3978
rect -7731 2107 -7615 2113
rect -14886 2093 -14822 2099
rect -14886 1002 -14822 2029
rect -7731 2013 -7725 2107
rect -7621 2013 -7615 2107
rect -5486 2042 -5358 2224
rect -7725 1595 -7621 2013
rect -7725 1539 -7696 1595
rect -7640 1539 -7621 1595
rect -14886 946 -14882 1002
rect -14826 946 -14822 1002
rect -14886 942 -14822 946
rect -13792 1006 -13728 1015
rect -14882 937 -14826 942
rect -13792 -614 -13728 942
rect -9252 -465 -9124 -456
rect -13792 -670 -13788 -614
rect -13732 -670 -13728 -614
rect -13792 -674 -13728 -670
rect -11294 -610 -11230 -601
rect -13788 -679 -13732 -674
rect -16333 -772 -16273 -763
rect -11470 -772 -11414 -765
rect -16333 -841 -16273 -832
rect -11472 -774 -11412 -772
rect -11472 -830 -11470 -774
rect -11414 -830 -11412 -774
rect -11648 -900 -11584 -891
rect -11648 -1490 -11584 -964
rect -11653 -1546 -11644 -1490
rect -11588 -1546 -11579 -1490
rect -11648 -1550 -11584 -1546
rect -11472 -1661 -11412 -830
rect -11476 -1670 -11412 -1661
rect -11420 -1726 -11412 -1670
rect -11476 -1735 -11412 -1726
rect -11294 -1841 -11230 -674
rect -11294 -1897 -11292 -1841
rect -11236 -1897 -11230 -1841
rect -11294 -1909 -11230 -1897
rect -9252 -1704 -9124 -593
rect -9252 -1756 -9246 -1704
rect -9130 -1756 -9124 -1704
rect -15351 -2196 -15287 -2068
rect -17666 -2734 -17657 -2678
rect -17601 -2734 -17592 -2678
rect -17661 -2738 -17597 -2734
rect -13162 -2745 -13084 -2709
rect -13162 -7524 -13098 -2745
rect -9252 -3438 -9124 -1756
rect -9252 -3490 -9246 -3438
rect -9130 -3490 -9124 -3438
rect -9252 -4344 -9124 -3490
rect -9252 -4532 -9246 -4344
rect -9130 -4532 -9124 -4344
rect -9252 -4538 -9124 -4532
rect -9052 -1430 -8924 -712
rect -9052 -1668 -9046 -1430
rect -8930 -1668 -8924 -1430
rect -9052 -3164 -8924 -1668
rect -9052 -3402 -9046 -3164
rect -8930 -3402 -8924 -3164
rect -9052 -4600 -8924 -3402
rect -9052 -4788 -9046 -4600
rect -8930 -4788 -8924 -4600
rect -9052 -4794 -8924 -4788
rect -8852 -718 -8724 -712
rect -8852 -854 -8846 -718
rect -8730 -854 -8724 -718
rect -8852 -2244 -8724 -854
rect -8047 -1933 -7983 -1927
rect -8047 -2049 -8041 -1933
rect -7989 -2049 -7983 -1933
rect -8047 -2119 -7983 -2049
rect -8852 -2588 -8846 -2244
rect -8730 -2588 -8724 -2244
rect -8852 -3978 -8724 -2588
rect -8047 -3667 -7983 -3661
rect -8047 -3783 -8041 -3667
rect -7989 -3783 -7983 -3667
rect -8047 -3853 -7983 -3783
rect -8852 -4114 -8846 -3978
rect -8730 -4114 -8724 -3978
rect -13162 -7580 -13158 -7524
rect -13102 -7580 -13098 -7524
rect -13162 -7584 -13098 -7580
rect -13158 -7589 -13102 -7584
rect -18588 -8100 -18586 -8044
rect -18530 -8100 -18528 -8044
rect -18588 -8102 -18528 -8100
rect -18586 -8109 -18530 -8102
rect -27806 -10796 -27800 -10519
rect -27412 -10796 -27406 -10519
rect -27806 -10802 -27406 -10796
rect -28262 -11096 -28256 -10858
rect -27868 -11096 -27862 -10858
rect -28262 -11102 -27862 -11096
rect -8852 -16902 -8724 -4114
rect -8318 -9078 -8224 -9074
rect -7725 -9078 -7621 1539
rect -5486 1883 -5478 2042
rect -5364 1883 -5358 2042
rect -5486 706 -5358 1883
rect -5486 630 -5477 706
rect -5370 630 -5358 706
rect -5486 -465 -5358 630
rect -5486 -599 -5358 -593
rect -5286 1397 -5158 2224
rect -4639 1604 -4583 1703
rect -4641 1595 -4583 1604
rect -4585 1539 -4583 1595
rect -4641 1530 -4583 1539
rect -4639 1472 -4583 1530
rect -5286 1240 -5277 1397
rect -5167 1240 -5158 1397
rect -5286 167 -5158 1240
rect -4230 1179 -4174 1186
rect -4232 1177 -4172 1179
rect -4232 1121 -4230 1177
rect -4174 1121 -4172 1177
rect -4232 896 -4172 1121
rect -4696 894 -4636 896
rect -4703 838 -4694 894
rect -4638 838 -4629 894
rect -4696 395 -4636 838
rect -4232 827 -4172 836
rect -3178 496 -3111 508
rect -3178 387 -3173 496
rect -4696 329 -4636 335
rect -3179 331 -3173 387
rect -3178 241 -3173 331
rect -3117 387 -3111 496
rect -3117 331 -2990 387
rect -3117 241 -3111 331
rect -3178 229 -3111 241
rect -5286 83 -5278 167
rect -5166 83 -5158 167
rect -5286 -732 -5158 83
rect -5286 -866 -5158 -860
rect -6515 -1201 -6451 -1195
rect -6515 -1317 -6509 -1201
rect -6457 -1317 -6451 -1201
rect -6515 -2796 -6451 -1317
rect -4403 -1201 -4339 -1195
rect -4403 -1317 -4397 -1201
rect -4345 -1317 -4339 -1201
rect -5935 -1933 -5871 -1927
rect -5935 -2049 -5929 -1933
rect -5877 -2049 -5871 -1933
rect -5935 -2119 -5871 -2049
rect -4403 -2767 -4339 -1317
rect -2291 -1201 -2227 -1195
rect -2291 -1317 -2285 -1201
rect -2233 -1317 -2227 -1201
rect -3823 -1933 -3759 -1927
rect -3823 -2049 -3817 -1933
rect -3765 -2049 -3759 -1933
rect -3823 -2119 -3759 -2049
rect -2291 -2745 -2227 -1317
rect -179 -1201 -115 -1195
rect -179 -1317 -173 -1201
rect -121 -1317 -115 -1201
rect -1711 -1933 -1647 -1927
rect -1711 -2049 -1705 -1933
rect -1653 -2049 -1647 -1933
rect -1711 -2119 -1647 -2049
rect -179 -2724 -115 -1317
rect 1933 -1201 1997 -1195
rect 1933 -1317 1939 -1201
rect 1991 -1317 1997 -1201
rect 401 -1933 465 -1927
rect 401 -2049 407 -1933
rect 459 -2049 465 -1933
rect 401 -2119 465 -2049
rect -6515 -2860 -6341 -2796
rect -4403 -2831 -4223 -2767
rect -2291 -2809 -2111 -2745
rect -179 -2788 44 -2724
rect -6515 -2935 -6451 -2929
rect -6515 -3051 -6509 -2935
rect -6457 -3051 -6451 -2935
rect -6515 -7297 -6451 -3051
rect -6405 -7158 -6341 -2860
rect -4403 -2935 -4339 -2929
rect -4403 -3051 -4397 -2935
rect -4345 -3051 -4339 -2935
rect -4403 -3489 -4339 -3051
rect -4287 -3470 -4223 -2831
rect -2291 -2935 -2227 -2929
rect -2291 -3051 -2285 -2935
rect -2233 -3051 -2227 -2935
rect -4403 -3529 -4338 -3489
rect -4287 -3519 -4222 -3470
rect -5935 -3667 -5871 -3661
rect -5935 -3783 -5929 -3667
rect -5877 -3783 -5871 -3667
rect -4402 -3702 -4338 -3529
rect -4286 -3569 -4222 -3519
rect -4286 -3625 -4282 -3569
rect -4226 -3625 -4222 -3569
rect -4286 -3629 -4222 -3625
rect -2618 -3565 -2554 -3556
rect -4282 -3634 -4226 -3629
rect -4402 -3758 -4398 -3702
rect -4342 -3758 -4338 -3702
rect -4402 -3762 -4338 -3758
rect -3823 -3667 -3759 -3661
rect -4398 -3767 -4342 -3762
rect -5935 -3853 -5871 -3783
rect -3823 -3783 -3817 -3667
rect -3765 -3783 -3759 -3667
rect -3823 -3853 -3759 -3783
rect -3146 -3698 -3082 -3689
rect -3666 -7152 -3610 -7147
rect -6405 -7231 -6341 -7222
rect -3670 -7156 -3606 -7152
rect -3670 -7212 -3666 -7156
rect -3610 -7212 -3606 -7156
rect -6515 -7370 -6451 -7361
rect -4212 -7302 -4156 -7293
rect -4212 -7367 -4156 -7358
rect -3670 -7371 -3606 -7212
rect -3146 -7382 -3082 -3762
rect -2618 -7374 -2554 -3629
rect -2291 -4510 -2227 -3051
rect -2175 -4344 -2111 -2809
rect -179 -2935 -115 -2929
rect -179 -3051 -173 -2935
rect -121 -3051 -115 -2935
rect -1711 -3667 -1647 -3661
rect -1711 -3783 -1705 -3667
rect -1653 -3783 -1647 -3667
rect -1711 -3853 -1647 -3783
rect -2175 -4417 -2111 -4408
rect -1533 -4344 -1469 -4335
rect -2291 -4583 -2227 -4574
rect -2083 -4511 -2019 -4502
rect -2083 -7374 -2019 -4575
rect -1533 -7374 -1469 -4408
rect -1003 -4826 -934 -4817
rect -1003 -7367 -934 -4895
rect -179 -4830 -115 -3051
rect -179 -4889 -173 -4830
rect -117 -4889 -115 -4830
rect -179 -4899 -115 -4889
rect -20 -4872 44 -2788
rect 1933 -2782 1997 -1317
rect 4045 -1201 4109 -1195
rect 4045 -1317 4051 -1201
rect 4103 -1317 4109 -1201
rect 2513 -1933 2577 -1927
rect 2513 -2049 2519 -1933
rect 2571 -2049 2577 -1933
rect 2513 -2119 2577 -2049
rect 4045 -2778 4109 -1317
rect 6157 -1201 6221 -1195
rect 6157 -1317 6163 -1201
rect 6215 -1317 6221 -1201
rect 4625 -1933 4689 -1927
rect 4625 -2049 4631 -1933
rect 4683 -2049 4689 -1933
rect 4625 -2119 4689 -2049
rect 6157 -2771 6221 -1317
rect 8269 -1201 8333 -1195
rect 8269 -1317 8275 -1201
rect 8327 -1317 8333 -1201
rect 6737 -1933 6801 -1927
rect 6737 -2049 6743 -1933
rect 6795 -2049 6801 -1933
rect 6737 -2119 6801 -2049
rect 8269 -2742 8333 -1317
rect 10381 -1201 10445 -1195
rect 10381 -1317 10387 -1201
rect 10439 -1317 10445 -1201
rect 10381 -1486 10445 -1317
rect 10381 -1559 10445 -1550
rect 10636 -1324 10696 -1318
rect 10636 -1670 10696 -1384
rect 10629 -1726 10638 -1670
rect 10694 -1726 10703 -1670
rect 10636 -1728 10696 -1726
rect 11174 -1837 11250 -1831
rect 11174 -1901 11180 -1837
rect 11244 -1901 11250 -1837
rect 11174 -1907 11250 -1901
rect 8849 -1933 8913 -1927
rect 8849 -2049 8855 -1933
rect 8907 -2049 8913 -1933
rect 8849 -2119 8913 -2049
rect 1933 -2846 2149 -2782
rect 4045 -2842 4247 -2778
rect 6157 -2835 6367 -2771
rect 8269 -2806 8480 -2742
rect 1933 -2935 1997 -2929
rect 1933 -3051 1939 -2935
rect 1991 -3051 1997 -2935
rect 401 -3667 465 -3661
rect 401 -3783 407 -3667
rect 459 -3783 465 -3667
rect 401 -3853 465 -3783
rect 1076 -3859 1132 -3854
rect 1933 -3859 1997 -3051
rect 1072 -3863 1136 -3859
rect 1072 -3919 1076 -3863
rect 1132 -3919 1136 -3863
rect -20 -4899 47 -4872
rect -479 -5097 -470 -5033
rect -406 -5097 -397 -5033
rect -17 -5037 47 -4899
rect -17 -5093 -13 -5037
rect 43 -5093 47 -5037
rect -17 -5097 47 -5093
rect -470 -7382 -406 -5097
rect -13 -5102 43 -5097
rect 72 -5202 136 -5193
rect 1072 -5206 1136 -3919
rect 1933 -3932 1997 -3923
rect 1597 -3997 1653 -3992
rect 2085 -3997 2149 -2846
rect 4045 -2935 4109 -2929
rect 4045 -3051 4051 -2935
rect 4103 -3051 4109 -2935
rect 2513 -3667 2577 -3661
rect 2513 -3783 2519 -3667
rect 2571 -3783 2577 -3667
rect 2513 -3853 2577 -3783
rect 1593 -4001 1657 -3997
rect 1593 -4057 1597 -4001
rect 1653 -4057 1657 -4001
rect 1593 -4872 1657 -4057
rect 2085 -4070 2149 -4061
rect 2140 -4157 2196 -4152
rect 4045 -4157 4109 -3051
rect 2136 -4161 2200 -4157
rect 2136 -4217 2140 -4161
rect 2196 -4217 2200 -4161
rect 2136 -4830 2200 -4217
rect 4045 -4230 4109 -4221
rect 2669 -4311 2725 -4306
rect 4183 -4311 4247 -2842
rect 6157 -2935 6221 -2929
rect 6157 -3051 6163 -2935
rect 6215 -3051 6221 -2935
rect 4625 -3667 4689 -3661
rect 4625 -3783 4631 -3667
rect 4683 -3783 4689 -3667
rect 4625 -3853 4689 -3783
rect 2665 -4315 2729 -4311
rect 2665 -4371 2669 -4315
rect 2725 -4371 2729 -4315
rect 1593 -4899 1658 -4872
rect 2136 -4899 2201 -4830
rect 1072 -5262 1076 -5206
rect 1132 -5262 1136 -5206
rect 1072 -5266 1136 -5262
rect 72 -7374 136 -5266
rect 1076 -5271 1132 -5266
rect 593 -5367 657 -5358
rect 1594 -5371 1658 -4899
rect 1594 -5427 1598 -5371
rect 1654 -5427 1658 -5371
rect 1594 -5431 1658 -5427
rect 593 -7367 657 -5431
rect 1598 -5436 1654 -5431
rect 1136 -5543 1200 -5534
rect 2137 -5547 2201 -4899
rect 2137 -5603 2141 -5547
rect 2197 -5603 2201 -5547
rect 2137 -5607 2201 -5603
rect 1136 -7332 1200 -5607
rect 2141 -5612 2197 -5607
rect 1665 -5732 1729 -5723
rect 2665 -5736 2729 -4371
rect 4183 -4384 4247 -4375
rect 3205 -4458 3261 -4453
rect 6157 -4458 6221 -3051
rect 3201 -4462 3265 -4458
rect 3201 -4518 3205 -4462
rect 3261 -4518 3265 -4462
rect 3201 -4802 3265 -4518
rect 6157 -4531 6221 -4522
rect 3747 -4612 3803 -4607
rect 6303 -4612 6367 -2835
rect 8269 -2935 8333 -2929
rect 8269 -3051 8275 -2935
rect 8327 -3051 8333 -2935
rect 6737 -3667 6801 -3661
rect 6737 -3783 6743 -3667
rect 6795 -3783 6801 -3667
rect 6737 -3853 6801 -3783
rect 3743 -4616 3807 -4612
rect 3743 -4672 3747 -4616
rect 3803 -4672 3807 -4616
rect 3743 -4791 3807 -4672
rect 6303 -4685 6367 -4676
rect 3201 -4899 3267 -4802
rect 3743 -4899 3810 -4791
rect 4275 -4796 4331 -4791
rect 8269 -4796 8333 -3051
rect 4271 -4800 4335 -4796
rect 4271 -4856 4275 -4800
rect 4331 -4856 4335 -4800
rect 4271 -4861 4335 -4856
rect 4271 -4899 4336 -4861
rect 8269 -4869 8333 -4860
rect 8416 -4850 8480 -2806
rect 10381 -2935 10445 -2929
rect 10381 -3051 10387 -2935
rect 10439 -3051 10445 -2935
rect 8849 -3667 8913 -3661
rect 8849 -3783 8855 -3667
rect 8907 -3783 8913 -3667
rect 8849 -3853 8913 -3783
rect 10381 -4841 10445 -3051
rect 8416 -4899 8481 -4850
rect 2665 -5792 2669 -5736
rect 2725 -5792 2729 -5736
rect 2665 -5796 2729 -5792
rect 1665 -7375 1729 -5796
rect 2669 -5801 2725 -5796
rect 2201 -5925 2265 -5916
rect 3203 -5929 3267 -4899
rect 3203 -5985 3207 -5929
rect 3263 -5985 3267 -5929
rect 3203 -5989 3267 -5985
rect 2201 -7382 2265 -5989
rect 3207 -5994 3263 -5989
rect 2743 -6094 2807 -6085
rect 3746 -6098 3810 -4899
rect 3746 -6154 3750 -6098
rect 3806 -6154 3810 -6098
rect 3746 -6158 3810 -6154
rect 2743 -7390 2807 -6158
rect 3750 -6163 3806 -6158
rect 3271 -6270 3335 -6261
rect 4272 -6274 4336 -4899
rect 4272 -6330 4276 -6274
rect 4332 -6330 4336 -6274
rect 4272 -6334 4336 -6330
rect 4424 -4984 4488 -4975
rect 8417 -4988 8481 -4899
rect 8417 -5044 8421 -4988
rect 8477 -5044 8481 -4988
rect 8417 -5048 8481 -5044
rect 10380 -4899 10445 -4841
rect 3271 -7368 3335 -6334
rect 4276 -6339 4332 -6334
rect 3801 -6421 3865 -6412
rect 4424 -6425 4488 -5048
rect 8421 -5053 8477 -5048
rect 4424 -6481 4428 -6425
rect 4484 -6481 4488 -6425
rect 4424 -6485 4488 -6481
rect 4571 -5188 4635 -5179
rect 10380 -5192 10444 -4899
rect 10380 -5248 10384 -5192
rect 10440 -5248 10444 -5192
rect 10380 -5252 10444 -5248
rect 3801 -7368 3865 -6485
rect 4428 -6490 4484 -6485
rect -5084 -7520 -5028 -7515
rect -5088 -7524 -5024 -7520
rect -5088 -7580 -5084 -7524
rect -5028 -7580 -5024 -7524
rect -5088 -8780 -5024 -7580
rect 4571 -7524 4635 -5252
rect 10384 -5257 10440 -5252
rect 4571 -7580 4575 -7524
rect 4631 -7580 4635 -7524
rect 4571 -7584 4635 -7580
rect 4575 -7589 4631 -7584
rect -4390 -8042 -4330 -8033
rect -4390 -8904 -4330 -8102
rect -4390 -8960 -4388 -8904
rect -4332 -8960 -4330 -8904
rect -4390 -8962 -4330 -8960
rect -4388 -8969 -4332 -8962
rect -8323 -9083 -8219 -9078
rect -8323 -9177 -8318 -9083
rect -8224 -9177 -8219 -9083
rect -8323 -16884 -8219 -9177
rect -7725 -9191 -7621 -9182
rect -7484 -9963 -7380 -9815
rect -5082 -10830 -4381 -10824
rect -5082 -11018 -5076 -10830
rect -4893 -11018 -4575 -10830
rect -4387 -11018 -4381 -10830
rect -5082 -11024 -4381 -11018
rect -8323 -16997 -8219 -16988
rect -8852 -17039 -8724 -17030
<< via2 >>
rect -29004 10118 -28866 10256
rect -27929 10119 -27868 10255
rect -29931 -1371 -29793 -1233
rect -19249 7687 -19185 7751
rect -27035 7091 -26979 7147
rect -27478 6676 -27412 6812
rect -27478 2178 -27412 2314
rect -17661 7087 -17597 7151
rect -18588 5454 -18528 5514
rect -18293 5250 -18229 5314
rect -15146 6807 -15090 6809
rect -15146 6681 -15144 6807
rect -15144 6681 -15092 6807
rect -15092 6681 -15090 6807
rect -15146 6679 -15090 6681
rect -4129 4678 -3999 4680
rect -4129 4552 -4127 4678
rect -4127 4552 -4001 4678
rect -4001 4552 -3999 4678
rect -4129 4550 -3999 4552
rect -3915 4604 -3859 4606
rect -3915 4552 -3913 4604
rect -3913 4552 -3861 4604
rect -3861 4552 -3859 4604
rect -3915 4550 -3859 4552
rect -3780 4678 -3724 4680
rect -3780 4552 -3778 4678
rect -3778 4552 -3726 4678
rect -3726 4552 -3724 4678
rect -3780 4550 -3724 4552
rect -4613 4302 -4483 4432
rect -4398 4302 -4342 4358
rect -4264 4302 -4208 4432
rect -4129 4430 -3999 4432
rect -4129 4304 -4127 4430
rect -4127 4304 -4001 4430
rect -4001 4304 -3999 4430
rect -4129 4302 -3999 4304
rect -3915 4356 -3859 4358
rect -3915 4304 -3913 4356
rect -3913 4304 -3861 4356
rect -3861 4304 -3859 4356
rect -3915 4302 -3859 4304
rect -3780 4430 -3724 4432
rect -3780 4304 -3778 4430
rect -3778 4304 -3726 4430
rect -3726 4304 -3724 4430
rect -3780 4302 -3724 4304
rect -4255 4022 -4125 4078
rect -3771 4032 -3641 4034
rect -3771 3980 -3769 4032
rect -3769 3980 -3643 4032
rect -3643 3980 -3641 4032
rect -3771 3978 -3641 3980
rect -7696 1539 -7640 1595
rect -14882 946 -14826 1002
rect -13792 942 -13728 1006
rect -13788 -670 -13732 -614
rect -11294 -674 -11230 -610
rect -16333 -832 -16273 -772
rect -11470 -830 -11414 -774
rect -11648 -964 -11584 -900
rect -11644 -1546 -11588 -1490
rect -11476 -1726 -11420 -1670
rect -11292 -1897 -11236 -1841
rect -17657 -2734 -17601 -2678
rect -13158 -7580 -13102 -7524
rect -18586 -8100 -18530 -8044
rect -4641 1539 -4585 1595
rect -4230 1121 -4174 1177
rect -4694 838 -4638 894
rect -4232 836 -4172 896
rect -4282 -3625 -4226 -3569
rect -2618 -3629 -2554 -3565
rect -4398 -3758 -4342 -3702
rect -3146 -3762 -3082 -3698
rect -6405 -7222 -6341 -7158
rect -3666 -7212 -3610 -7156
rect -6515 -7361 -6451 -7297
rect -4212 -7358 -4156 -7302
rect -2175 -4408 -2111 -4344
rect -1533 -4408 -1469 -4344
rect -2291 -4574 -2227 -4510
rect -2083 -4575 -2019 -4511
rect -1003 -4895 -934 -4826
rect -173 -4889 -117 -4830
rect 10381 -1550 10445 -1486
rect 10638 -1726 10694 -1670
rect 11184 -1897 11240 -1841
rect 1076 -3919 1132 -3863
rect -470 -5097 -406 -5033
rect -13 -5093 43 -5037
rect 72 -5266 136 -5202
rect 1933 -3923 1997 -3859
rect 1597 -4057 1653 -4001
rect 2085 -4061 2149 -3997
rect 2140 -4217 2196 -4161
rect 4045 -4221 4109 -4157
rect 2669 -4371 2725 -4315
rect 1076 -5262 1132 -5206
rect 593 -5431 657 -5367
rect 1598 -5427 1654 -5371
rect 1136 -5607 1200 -5543
rect 2141 -5603 2197 -5547
rect 1665 -5796 1729 -5732
rect 4183 -4375 4247 -4311
rect 3205 -4518 3261 -4462
rect 6157 -4522 6221 -4458
rect 3747 -4672 3803 -4616
rect 6303 -4676 6367 -4612
rect 4275 -4856 4331 -4800
rect 8269 -4860 8333 -4796
rect 2669 -5792 2725 -5736
rect 2201 -5989 2265 -5925
rect 3207 -5985 3263 -5929
rect 2743 -6158 2807 -6094
rect 3750 -6154 3806 -6098
rect 3271 -6334 3335 -6270
rect 4276 -6330 4332 -6274
rect 4424 -5048 4488 -4984
rect 8421 -5044 8477 -4988
rect 3801 -6485 3865 -6421
rect 4428 -6481 4484 -6425
rect 4571 -5252 4635 -5188
rect 10384 -5248 10440 -5192
rect -5084 -7580 -5028 -7524
rect 4575 -7580 4631 -7524
rect -4390 -8102 -4330 -8042
rect -4388 -8960 -4332 -8904
rect -8852 -17030 -8724 -16902
rect -8318 -9177 -8224 -9083
rect -7725 -9182 -7621 -9078
rect -8323 -16988 -8219 -16884
<< metal3 >>
rect -29009 10256 -27136 10261
rect -29009 10118 -29004 10256
rect -28866 10255 -27136 10256
rect -28866 10119 -27929 10255
rect -27868 10119 -27136 10255
rect -28866 10118 -27136 10119
rect -29009 10113 -27136 10118
rect -27218 7751 -19180 7756
rect -27218 7687 -19249 7751
rect -19185 7687 -19180 7751
rect -27218 7682 -19180 7687
rect -27040 7151 -26974 7152
rect -17666 7151 -17592 7156
rect -27040 7147 -17661 7151
rect -27040 7091 -27035 7147
rect -26979 7091 -17661 7147
rect -27040 7087 -17661 7091
rect -17597 7087 -17592 7151
rect -27040 7086 -26974 7087
rect -17666 7082 -17592 7087
rect -27484 6812 -27166 6818
rect -27484 6676 -27478 6812
rect -27412 6676 -27166 6812
rect -27484 6670 -27166 6676
rect -15503 6809 -15081 6818
rect -15503 6679 -15146 6809
rect -15090 6679 -15081 6809
rect -15503 6670 -15081 6679
rect -18593 5514 -18523 5519
rect -18593 5454 -18588 5514
rect -18528 5454 -18523 5514
rect -18593 5449 -18523 5454
rect -18298 5314 -18224 5319
rect -18298 5250 -18293 5314
rect -18229 5250 -18224 5314
rect -18298 5245 -18224 5250
rect -4138 4680 -3990 4689
rect -4138 4550 -4129 4680
rect -3999 4550 -3990 4680
rect -3789 4680 -3715 4689
rect -4138 4541 -3990 4550
rect -3924 4606 -3850 4615
rect -3924 4550 -3915 4606
rect -3859 4550 -3850 4606
rect -3924 4541 -3850 4550
rect -3789 4550 -3780 4680
rect -3724 4550 -3715 4680
rect -3789 4541 -3715 4550
rect -4622 4432 -4474 4441
rect -4622 4302 -4613 4432
rect -4483 4302 -4474 4432
rect -4273 4432 -4199 4441
rect -4622 4293 -4474 4302
rect -4407 4358 -4333 4367
rect -4407 4302 -4398 4358
rect -4342 4302 -4333 4358
rect -4407 4293 -4333 4302
rect -4273 4302 -4264 4432
rect -4208 4302 -4199 4432
rect -4273 4293 -4199 4302
rect -4138 4432 -3990 4441
rect -4138 4302 -4129 4432
rect -3999 4302 -3990 4432
rect -3789 4432 -3715 4441
rect -4138 4293 -3990 4302
rect -3924 4358 -3850 4367
rect -3924 4302 -3915 4358
rect -3859 4302 -3850 4358
rect -3924 4293 -3850 4302
rect -3789 4302 -3780 4432
rect -3724 4302 -3715 4432
rect -3789 4293 -3715 4302
rect -4264 4078 -4116 4087
rect -4264 4022 -4255 4078
rect -4125 4022 -4116 4078
rect -4264 4013 -4116 4022
rect -3780 4034 -3632 4043
rect -3780 3978 -3771 4034
rect -3641 3978 -3632 4034
rect -3780 3969 -3632 3978
rect -27484 2314 -26420 2320
rect -27484 2178 -27478 2314
rect -27412 2178 -26420 2314
rect -27484 2172 -26420 2178
rect -7701 1597 -7635 1600
rect -4646 1597 -4580 1600
rect -7701 1595 -4580 1597
rect -7701 1539 -7696 1595
rect -7640 1539 -4641 1595
rect -4585 1539 -4580 1595
rect -7701 1537 -4580 1539
rect -7701 1534 -7635 1537
rect -4646 1534 -4580 1537
rect -4235 1179 -4169 1182
rect -4235 1177 -3974 1179
rect -4235 1121 -4230 1177
rect -4174 1121 -3974 1177
rect -4235 1119 -3974 1121
rect -4235 1116 -4169 1119
rect -14887 1006 -14821 1007
rect -13797 1006 -13723 1011
rect -14887 1002 -13792 1006
rect -14887 946 -14882 1002
rect -14826 946 -13792 1002
rect -14887 942 -13792 946
rect -13728 942 -13723 1006
rect -14887 941 -14821 942
rect -13797 937 -13723 942
rect -4699 896 -4633 899
rect -4237 896 -4167 901
rect -4699 894 -4232 896
rect -4699 838 -4694 894
rect -4638 838 -4232 894
rect -4699 836 -4232 838
rect -4172 836 -4167 896
rect -4699 833 -4633 836
rect -4237 831 -4167 836
rect -13793 -610 -13727 -609
rect -11299 -610 -11225 -605
rect -13793 -614 -11294 -610
rect -13793 -670 -13788 -614
rect -13732 -670 -11294 -614
rect -13793 -674 -11294 -670
rect -11230 -674 -11225 -610
rect -13793 -675 -13727 -674
rect -11299 -679 -11225 -674
rect -16338 -772 -16268 -767
rect -11475 -772 -11409 -769
rect -16338 -832 -16333 -772
rect -16273 -774 -11409 -772
rect -16273 -830 -11470 -774
rect -11414 -830 -11409 -774
rect -16273 -832 -11409 -830
rect -16338 -837 -16268 -832
rect -11475 -835 -11409 -832
rect -11653 -900 -11579 -895
rect -11771 -964 -11648 -900
rect -11584 -964 -11579 -900
rect -11653 -969 -11579 -964
rect -29936 -1233 -26949 -1228
rect -29936 -1371 -29931 -1233
rect -29793 -1371 -26949 -1233
rect -29936 -1376 -26949 -1371
rect -11649 -1486 -11583 -1485
rect 10376 -1486 10450 -1481
rect -11649 -1490 10381 -1486
rect -11649 -1546 -11644 -1490
rect -11588 -1546 10381 -1490
rect -11649 -1550 10381 -1546
rect 10445 -1550 10450 -1486
rect -11649 -1551 -11583 -1550
rect 10376 -1555 10450 -1550
rect -11481 -1668 -11415 -1665
rect 10633 -1668 10699 -1665
rect -11481 -1670 10699 -1668
rect -11481 -1726 -11476 -1670
rect -11420 -1726 10638 -1670
rect 10694 -1726 10699 -1670
rect -11481 -1728 10699 -1726
rect -11481 -1731 -11415 -1728
rect 10633 -1731 10699 -1728
rect -11297 -1837 -11231 -1836
rect 11174 -1837 11250 -1831
rect -11297 -1841 11250 -1837
rect -11297 -1897 -11292 -1841
rect -11236 -1897 11184 -1841
rect 11240 -1897 11250 -1841
rect -11297 -1901 11250 -1897
rect -11297 -1902 -11231 -1901
rect 11174 -1907 11250 -1901
rect -17662 -2674 -17596 -2673
rect -17662 -2678 -15348 -2674
rect -17662 -2734 -17657 -2678
rect -17601 -2734 -15348 -2678
rect -17662 -2738 -15348 -2734
rect -17662 -2739 -17596 -2738
rect -15414 -2793 -15348 -2738
rect -15414 -2858 -15412 -2793
rect -4287 -3565 -4221 -3564
rect -2623 -3565 -2549 -3560
rect -4287 -3569 -2618 -3565
rect -4287 -3625 -4282 -3569
rect -4226 -3625 -2618 -3569
rect -4287 -3629 -2618 -3625
rect -2554 -3629 -2549 -3565
rect -4287 -3630 -4221 -3629
rect -2623 -3634 -2549 -3629
rect -4403 -3698 -4337 -3697
rect -3151 -3698 -3077 -3693
rect -4403 -3702 -3146 -3698
rect -4403 -3758 -4398 -3702
rect -4342 -3758 -3146 -3702
rect -4403 -3762 -3146 -3758
rect -3082 -3762 -3077 -3698
rect -4403 -3763 -4337 -3762
rect -3151 -3767 -3077 -3762
rect 1071 -3859 1137 -3858
rect 1928 -3859 2002 -3854
rect 1071 -3863 1933 -3859
rect 1071 -3919 1076 -3863
rect 1132 -3919 1933 -3863
rect 1071 -3923 1933 -3919
rect 1997 -3923 2002 -3859
rect 1071 -3924 1137 -3923
rect 1928 -3928 2002 -3923
rect 1592 -3997 1658 -3996
rect 2080 -3997 2154 -3992
rect 1592 -4001 2085 -3997
rect 1592 -4057 1597 -4001
rect 1653 -4057 2085 -4001
rect 1592 -4061 2085 -4057
rect 2149 -4061 2154 -3997
rect 1592 -4062 1658 -4061
rect 2080 -4066 2154 -4061
rect 2135 -4157 2201 -4156
rect 4040 -4157 4114 -4152
rect 2135 -4161 4045 -4157
rect 2135 -4217 2140 -4161
rect 2196 -4217 4045 -4161
rect 2135 -4221 4045 -4217
rect 4109 -4221 4114 -4157
rect 2135 -4222 2201 -4221
rect 4040 -4226 4114 -4221
rect 2664 -4311 2730 -4310
rect 4178 -4311 4252 -4306
rect 2664 -4315 4183 -4311
rect -2180 -4344 -2106 -4339
rect -1538 -4344 -1464 -4339
rect -2180 -4408 -2175 -4344
rect -2111 -4408 -1533 -4344
rect -1469 -4408 -1464 -4344
rect 2664 -4371 2669 -4315
rect 2725 -4371 4183 -4315
rect 2664 -4375 4183 -4371
rect 4247 -4375 4252 -4311
rect 2664 -4376 2730 -4375
rect 4178 -4380 4252 -4375
rect -2180 -4413 -2106 -4408
rect -1538 -4413 -1464 -4408
rect 3200 -4458 3266 -4457
rect 6152 -4458 6226 -4453
rect 3200 -4462 6157 -4458
rect -2296 -4510 -2222 -4505
rect -2088 -4510 -2014 -4506
rect -2296 -4574 -2291 -4510
rect -2227 -4511 -2014 -4510
rect -2227 -4574 -2083 -4511
rect -2296 -4579 -2222 -4574
rect -2088 -4575 -2083 -4574
rect -2019 -4575 -2014 -4511
rect 3200 -4518 3205 -4462
rect 3261 -4518 6157 -4462
rect 3200 -4522 6157 -4518
rect 6221 -4522 6226 -4458
rect 3200 -4523 3266 -4522
rect 6152 -4527 6226 -4522
rect -2088 -4580 -2014 -4575
rect 3742 -4612 3808 -4611
rect 6298 -4612 6372 -4607
rect 3742 -4616 6303 -4612
rect 3742 -4672 3747 -4616
rect 3803 -4672 6303 -4616
rect 3742 -4676 6303 -4672
rect 6367 -4676 6372 -4612
rect 3742 -4677 3808 -4676
rect 6298 -4681 6372 -4676
rect 4270 -4796 4336 -4795
rect 8264 -4796 8338 -4791
rect 4270 -4800 8269 -4796
rect -1008 -4825 -929 -4821
rect -1008 -4826 -112 -4825
rect -1008 -4895 -1003 -4826
rect -934 -4830 -112 -4826
rect -934 -4889 -173 -4830
rect -117 -4889 -112 -4830
rect 4270 -4856 4275 -4800
rect 4331 -4856 8269 -4800
rect 4270 -4860 8269 -4856
rect 8333 -4860 8338 -4796
rect 4270 -4861 4336 -4860
rect 8264 -4865 8338 -4860
rect -934 -4894 -112 -4889
rect -934 -4895 -929 -4894
rect -1008 -4900 -929 -4895
rect 4419 -4984 4493 -4979
rect 8416 -4984 8482 -4983
rect -475 -5033 -401 -5028
rect -18 -5033 48 -5032
rect -475 -5097 -470 -5033
rect -406 -5037 48 -5033
rect -406 -5093 -13 -5037
rect 43 -5093 48 -5037
rect 4419 -5048 4424 -4984
rect 4488 -4988 8482 -4984
rect 4488 -5044 8421 -4988
rect 8477 -5044 8482 -4988
rect 4488 -5048 8482 -5044
rect 4419 -5053 4493 -5048
rect 8416 -5049 8482 -5048
rect -406 -5097 48 -5093
rect -475 -5102 -401 -5097
rect -18 -5098 48 -5097
rect 4566 -5188 4640 -5183
rect 10379 -5188 10445 -5187
rect 67 -5202 141 -5197
rect 1071 -5202 1137 -5201
rect 67 -5266 72 -5202
rect 136 -5206 1137 -5202
rect 136 -5262 1076 -5206
rect 1132 -5262 1137 -5206
rect 4566 -5252 4571 -5188
rect 4635 -5192 10445 -5188
rect 4635 -5248 10384 -5192
rect 10440 -5248 10445 -5192
rect 4635 -5252 10445 -5248
rect 4566 -5257 4640 -5252
rect 10379 -5253 10445 -5252
rect 136 -5266 1137 -5262
rect 67 -5271 141 -5266
rect 1071 -5267 1137 -5266
rect 588 -5367 662 -5362
rect 1593 -5367 1659 -5366
rect 588 -5431 593 -5367
rect 657 -5371 1659 -5367
rect 657 -5427 1598 -5371
rect 1654 -5427 1659 -5371
rect 657 -5431 1659 -5427
rect 588 -5436 662 -5431
rect 1593 -5432 1659 -5431
rect 1131 -5543 1205 -5538
rect 2136 -5543 2202 -5542
rect 1131 -5607 1136 -5543
rect 1200 -5547 2202 -5543
rect 1200 -5603 2141 -5547
rect 2197 -5603 2202 -5547
rect 1200 -5607 2202 -5603
rect 1131 -5612 1205 -5607
rect 2136 -5608 2202 -5607
rect 1660 -5732 1734 -5727
rect 2664 -5732 2730 -5731
rect 1660 -5796 1665 -5732
rect 1729 -5736 2730 -5732
rect 1729 -5792 2669 -5736
rect 2725 -5792 2730 -5736
rect 1729 -5796 2730 -5792
rect 1660 -5801 1734 -5796
rect 2664 -5797 2730 -5796
rect 2196 -5925 2270 -5920
rect 3202 -5925 3268 -5924
rect 2196 -5989 2201 -5925
rect 2265 -5929 3268 -5925
rect 2265 -5985 3207 -5929
rect 3263 -5985 3268 -5929
rect 2265 -5989 3268 -5985
rect 2196 -5994 2270 -5989
rect 3202 -5990 3268 -5989
rect 2738 -6094 2812 -6089
rect 3745 -6094 3811 -6093
rect 2738 -6158 2743 -6094
rect 2807 -6098 3811 -6094
rect 2807 -6154 3750 -6098
rect 3806 -6154 3811 -6098
rect 2807 -6158 3811 -6154
rect 2738 -6163 2812 -6158
rect 3745 -6159 3811 -6158
rect 3266 -6270 3340 -6265
rect 4271 -6270 4337 -6269
rect 3266 -6334 3271 -6270
rect 3335 -6274 4337 -6270
rect 3335 -6330 4276 -6274
rect 4332 -6330 4337 -6274
rect 3335 -6334 4337 -6330
rect 3266 -6339 3340 -6334
rect 4271 -6335 4337 -6334
rect 3796 -6421 3870 -6416
rect 4423 -6421 4489 -6420
rect 3796 -6485 3801 -6421
rect 3865 -6425 4489 -6421
rect 3865 -6481 4428 -6425
rect 4484 -6481 4489 -6425
rect 3865 -6485 4489 -6481
rect 3796 -6490 3870 -6485
rect 4423 -6486 4489 -6485
rect -3671 -7152 -3605 -7151
rect -6410 -7156 -3605 -7152
rect -6410 -7158 -3666 -7156
rect -6410 -7222 -6405 -7158
rect -6341 -7212 -3666 -7158
rect -3610 -7212 -3605 -7156
rect -6341 -7216 -3605 -7212
rect -6341 -7222 -6336 -7216
rect -3671 -7217 -3605 -7216
rect -6410 -7227 -6336 -7222
rect -6520 -7297 -6446 -7292
rect -6520 -7361 -6515 -7297
rect -6451 -7298 -6446 -7297
rect -4217 -7298 -4151 -7297
rect -6451 -7302 -4151 -7298
rect -6451 -7358 -4212 -7302
rect -4156 -7358 -4151 -7302
rect -6451 -7361 -4151 -7358
rect -6520 -7362 -4151 -7361
rect -6520 -7366 -6446 -7362
rect -4217 -7363 -4151 -7362
rect -13163 -7520 -13097 -7519
rect -5089 -7520 -5023 -7519
rect 4570 -7520 4636 -7519
rect -13163 -7524 4636 -7520
rect -13163 -7580 -13158 -7524
rect -13102 -7580 -5084 -7524
rect -5028 -7580 4575 -7524
rect 4631 -7580 4636 -7524
rect -13163 -7584 4636 -7580
rect -13163 -7585 -13097 -7584
rect -5089 -7585 -5023 -7584
rect 4570 -7585 4636 -7584
rect -18591 -8042 -18525 -8039
rect -4395 -8042 -4325 -8037
rect -18591 -8044 -4390 -8042
rect -18591 -8100 -18586 -8044
rect -18530 -8100 -4390 -8044
rect -18591 -8102 -4390 -8100
rect -4330 -8102 -4325 -8042
rect -18591 -8105 -18525 -8102
rect -4395 -8107 -4325 -8102
rect -4393 -8902 -4327 -8899
rect -4393 -8904 -3729 -8902
rect -4393 -8960 -4388 -8904
rect -4332 -8960 -3729 -8904
rect -4393 -8962 -3729 -8960
rect 3724 -8962 3784 -8902
rect -4393 -8965 -4327 -8962
rect -7730 -9078 -7616 -9073
rect -8323 -9083 -7725 -9078
rect -8323 -9177 -8318 -9083
rect -8224 -9177 -7725 -9083
rect -8323 -9182 -7725 -9177
rect -7621 -9182 -7616 -9078
rect -7730 -9187 -7616 -9182
rect -8328 -16884 -8214 -16879
rect -6938 -16884 11081 -16882
rect -8863 -17035 -8857 -16897
rect -8729 -16902 -8719 -16897
rect -8724 -17030 -8719 -16902
rect -8328 -16988 -8323 -16884
rect -8219 -16986 11081 -16884
rect 11185 -16986 11191 -16882
rect -8219 -16988 -6884 -16986
rect -8328 -16993 -8214 -16988
rect -8729 -17035 -8719 -17030
<< via3 >>
rect -8857 -16902 -8729 -16897
rect -8857 -17030 -8852 -16902
rect -8852 -17030 -8729 -16902
rect 11081 -16986 11185 -16882
rect -8857 -17035 -8729 -17030
<< metal4 >>
rect 11080 -16882 11186 -16881
rect 11080 -16986 11081 -16882
rect 11185 -16986 11186 -16882
rect 11080 -16987 11186 -16986
rect 11081 -20941 11185 -16987
<< via4 >>
rect -8953 -16897 -8633 -16806
rect -8953 -17035 -8857 -16897
rect -8857 -17035 -8729 -16897
rect -8729 -17035 -8633 -16897
rect -8953 -17126 -8633 -17035
rect 10973 -21261 11293 -20941
<< metal5 >>
rect -8977 -16806 -8609 -16782
rect -8977 -17126 -8953 -16806
rect -8633 -17126 -8609 -16806
rect -8977 -17458 -8609 -17126
rect 10949 -20938 11317 -20917
rect 10345 -20941 11317 -20938
rect 10345 -21258 10973 -20941
rect 10949 -21261 10973 -21258
rect 11293 -21261 11317 -20941
rect 10949 -21285 11317 -21261
use comparator  comparator_0
timestamp 1712450145
transform 1 0 -26517 0 1 2397
box -811 -518 11035 7864
use ibias_gen  ibias_gen_0
timestamp 1712502012
transform 1 0 -27321 0 1 -10450
box -3279 -652 15828 11500
use rstring_mux  rstring_mux_0
timestamp 1712467038
transform 1 0 -16753 0 1 -15968
box -11632 -32 28451 9182
use schmitt_trigger  schmitt_trigger_0
timestamp 1712450145
transform 1 0 -4972 0 1 921
box -91 -52 2297 1163
use sky130_fd_pr__cap_mim_m3_2_LUWKLG  sky130_fd_pr__cap_mim_m3_2_LUWKLG_0
timestamp 1712463840
transform 0 -1 -8855 1 0 -20829
box -3349 -19200 3371 19200
use sky130_fd_pr__res_xhigh_po_1p41_DVQADA  sky130_fd_pr__res_xhigh_po_1p41_DVQADA_0
timestamp 1712352531
transform 1 0 -11267 0 1 5911
box -3898 -4082 3898 4082
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 -4929 0 1 125
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 -4469 0 1 125
box -38 -48 1510 592
use sky130_fd_sc_hvl__lsbufhv2lv_1  sky130_fd_sc_hvl__lsbufhv2lv_1_0
timestamp 1712419324
transform 1 0 10485 0 1 -2363
box -66 -43 1698 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 8 2112 0 1 1734
timestamp 1707688321
transform 1 0 -8523 0 1 -4097
box -66 -43 2178 1671
<< labels >>
flabel metal1 s -4580 -7558 -4580 -7558 0 FreeSans 1200 0 0 0 avss
port 20 nsew
flabel metal3 s 3724 -8962 3784 -8902 0 FreeSans 1200 0 0 0 vin
port 24 nsew
flabel metal2 -17531 753 -17531 753 0 FreeSans 1200 0 0 0 itest
port 25 nsew
flabel metal2 s -18241 -2814 -18241 -2814 0 FreeSans 1200 0 0 0 vbg_1v2
port 17 nsew
flabel metal2 -15287 -2068 -15287 -2068 0 FreeSans 1200 0 0 0 ibg_200n
port 26 nsew
flabel metal3 s 10400 -1728 10400 -1728 0 FreeSans 800 0 0 0 dcomp
flabel metal3 10912 -1837 10912 -1837 0 FreeSans 800 0 0 0 vl
flabel metal2 s 8849 -2119 8909 -2059 0 FreeSans 1200 0 0 0 isrc_sel
port 22 nsew
flabel metal2 s 8849 -3853 8909 -3793 0 FreeSans 1200 0 0 0 ena
port 18 nsew
flabel metal1 s -3836 -4436 -3836 -4436 0 FreeSans 1200 0 0 0 dvdd
port 21 nsew
flabel metal1 s -3836 -4646 -3836 -4646 0 FreeSans 1200 0 0 0 avdd
port 19 nsew
flabel metal2 s -8047 -2119 -8047 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[1]
port 15 nsew
flabel metal2 s -5935 -2119 -5935 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[3]
port 13 nsew
flabel metal2 s -3823 -2119 -3823 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[5]
port 11 nsew
flabel metal2 s -1711 -2119 -1711 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[7]
port 9 nsew
flabel metal2 s 401 -2119 401 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[9]
port 7 nsew
flabel metal2 s 2513 -2119 2513 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[11]
port 5 nsew
flabel metal2 s 4625 -2119 4625 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[13]
port 3 nsew
flabel metal2 s 6737 -2119 6737 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[15]
port 1 nsew
flabel metal2 s 6737 -3853 6737 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[14]
port 2 nsew
flabel metal2 s 4625 -3853 4625 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[12]
port 4 nsew
flabel metal2 s 2513 -3853 2513 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[10]
port 6 nsew
flabel metal2 s 401 -3853 401 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[8]
port 8 nsew
flabel metal2 s -1711 -3853 -1711 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[6]
port 10 nsew
flabel metal2 s -3823 -3853 -3823 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[4]
port 12 nsew
flabel metal2 s -5935 -3853 -5935 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[2]
port 14 nsew
flabel metal2 s -8047 -3853 -8047 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[0]
port 16 nsew
flabel metal2 -2990 331 -2990 331 0 FreeSans 1200 0 0 0 ovout
port 27 nsew
flabel metal2 -5158 -66 -5158 -66 0 FreeSans 1200 0 0 0 dvss
port 23 nsew
<< end >>
