magic
tech sky130A
magscale 1 2
timestamp 1712239005
<< metal4 >>
rect -10447 3039 -3749 3080
rect -10447 -3039 -4005 3039
rect -3769 -3039 -3749 3039
rect -10447 -3080 -3749 -3039
rect -3349 3039 3349 3080
rect -3349 -3039 3093 3039
rect 3329 -3039 3349 3039
rect -3349 -3080 3349 -3039
rect 3749 3039 10447 3080
rect 3749 -3039 10191 3039
rect 10427 -3039 10447 3039
rect 3749 -3080 10447 -3039
<< via4 >>
rect -4005 -3039 -3769 3039
rect 3093 -3039 3329 3039
rect 10191 -3039 10427 3039
<< mimcap2 >>
rect -10367 2960 -4367 3000
rect -10367 -2960 -10327 2960
rect -4407 -2960 -4367 2960
rect -10367 -3000 -4367 -2960
rect -3269 2960 2731 3000
rect -3269 -2960 -3229 2960
rect 2691 -2960 2731 2960
rect -3269 -3000 2731 -2960
rect 3829 2960 9829 3000
rect 3829 -2960 3869 2960
rect 9789 -2960 9829 2960
rect 3829 -3000 9829 -2960
<< mimcap2contact >>
rect -10327 -2960 -4407 2960
rect -3229 -2960 2691 2960
rect 3869 -2960 9789 2960
<< metal5 >>
rect -4047 3039 -3727 3081
rect -10351 2960 -4383 2984
rect -10351 -2960 -10327 2960
rect -4407 -2960 -4383 2960
rect -10351 -2984 -4383 -2960
rect -4047 -3039 -4005 3039
rect -3769 -3039 -3727 3039
rect 3051 3039 3371 3081
rect -3253 2960 2715 2984
rect -3253 -2960 -3229 2960
rect 2691 -2960 2715 2960
rect -3253 -2984 2715 -2960
rect -4047 -3081 -3727 -3039
rect 3051 -3039 3093 3039
rect 3329 -3039 3371 3039
rect 10149 3039 10469 3081
rect 3845 2960 9813 2984
rect 3845 -2960 3869 2960
rect 9789 -2960 9813 2960
rect 3845 -2984 9813 -2960
rect 3051 -3081 3371 -3039
rect 10149 -3039 10191 3039
rect 10427 -3039 10469 3039
rect 10149 -3081 10469 -3039
<< properties >>
string FIXED_BBOX 3749 -3080 9909 3080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 3 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
