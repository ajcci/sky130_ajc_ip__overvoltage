magic
tech sky130A
magscale 1 2
timestamp 1712463840
<< metal4 >>
rect -21094 3039 -14396 3080
rect -21094 -3039 -14652 3039
rect -14416 -3039 -14396 3039
rect -21094 -3080 -14396 -3039
rect -13996 3039 -7298 3080
rect -13996 -3039 -7554 3039
rect -7318 -3039 -7298 3039
rect -13996 -3080 -7298 -3039
rect -6898 3039 -200 3080
rect -6898 -3039 -456 3039
rect -220 -3039 -200 3039
rect -6898 -3080 -200 -3039
rect 200 3039 6898 3080
rect 200 -3039 6642 3039
rect 6878 -3039 6898 3039
rect 200 -3080 6898 -3039
rect 7298 3039 13996 3080
rect 7298 -3039 13740 3039
rect 13976 -3039 13996 3039
rect 7298 -3080 13996 -3039
rect 14396 3039 21094 3080
rect 14396 -3039 20838 3039
rect 21074 -3039 21094 3039
rect 14396 -3080 21094 -3039
<< via4 >>
rect -14652 -3039 -14416 3039
rect -7554 -3039 -7318 3039
rect -456 -3039 -220 3039
rect 6642 -3039 6878 3039
rect 13740 -3039 13976 3039
rect 20838 -3039 21074 3039
<< mimcap2 >>
rect -21014 2960 -15014 3000
rect -21014 -2960 -20974 2960
rect -15054 -2960 -15014 2960
rect -21014 -3000 -15014 -2960
rect -13916 2960 -7916 3000
rect -13916 -2960 -13876 2960
rect -7956 -2960 -7916 2960
rect -13916 -3000 -7916 -2960
rect -6818 2960 -818 3000
rect -6818 -2960 -6778 2960
rect -858 -2960 -818 2960
rect -6818 -3000 -818 -2960
rect 280 2960 6280 3000
rect 280 -2960 320 2960
rect 6240 -2960 6280 2960
rect 280 -3000 6280 -2960
rect 7378 2960 13378 3000
rect 7378 -2960 7418 2960
rect 13338 -2960 13378 2960
rect 7378 -3000 13378 -2960
rect 14476 2960 20476 3000
rect 14476 -2960 14516 2960
rect 20436 -2960 20476 2960
rect 14476 -3000 20476 -2960
<< mimcap2contact >>
rect -20974 -2960 -15054 2960
rect -13876 -2960 -7956 2960
rect -6778 -2960 -858 2960
rect 320 -2960 6240 2960
rect 7418 -2960 13338 2960
rect 14516 -2960 20436 2960
<< metal5 >>
rect -14694 3039 -14374 3081
rect -20998 2960 -15030 2984
rect -20998 -2960 -20974 2960
rect -15054 -2960 -15030 2960
rect -20998 -2984 -15030 -2960
rect -14694 -3039 -14652 3039
rect -14416 -3039 -14374 3039
rect -7596 3039 -7276 3081
rect -13900 2960 -7932 2984
rect -13900 -2960 -13876 2960
rect -7956 -2960 -7932 2960
rect -13900 -2984 -7932 -2960
rect -14694 -3081 -14374 -3039
rect -7596 -3039 -7554 3039
rect -7318 -3039 -7276 3039
rect -498 3039 -178 3081
rect -6802 2960 -834 2984
rect -6802 -2960 -6778 2960
rect -858 -2960 -834 2960
rect -6802 -2984 -834 -2960
rect -7596 -3081 -7276 -3039
rect -498 -3039 -456 3039
rect -220 -3039 -178 3039
rect 6600 3039 6920 3081
rect 296 2960 6264 2984
rect 296 -2960 320 2960
rect 6240 -2960 6264 2960
rect 296 -2984 6264 -2960
rect -498 -3081 -178 -3039
rect 6600 -3039 6642 3039
rect 6878 -3039 6920 3039
rect 13698 3039 14018 3081
rect 7394 2960 13362 2984
rect 7394 -2960 7418 2960
rect 13338 -2960 13362 2960
rect 7394 -2984 13362 -2960
rect 6600 -3081 6920 -3039
rect 13698 -3039 13740 3039
rect 13976 -3039 14018 3039
rect 20796 3039 21116 3081
rect 14492 2960 20460 2984
rect 14492 -2960 14516 2960
rect 20436 -2960 20460 2960
rect 14492 -2984 20460 -2960
rect 13698 -3081 14018 -3039
rect 20796 -3039 20838 3039
rect 21074 -3039 21116 3039
rect 20796 -3081 21116 -3039
<< properties >>
string FIXED_BBOX 14396 -3080 20556 3080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 6 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
