magic
tech sky130A
magscale 1 2
timestamp 1712450145
<< dnwell >>
rect -438 -438 10654 2526
<< nwell >>
rect -357 6707 -341 6741
rect -518 2320 10734 2606
rect -518 -232 -232 2320
rect 10448 -232 10734 2320
rect -518 -518 10734 -232
<< pwell >>
rect -386 4445 -322 4606
rect -515 4381 -322 4445
rect -515 3689 -451 4337
<< nsubdiff >>
rect -481 2549 10697 2569
rect -481 2515 -401 2549
rect 10617 2515 10697 2549
rect -481 2495 10697 2515
rect -481 2489 -407 2495
rect -481 -401 -461 2489
rect -427 -401 -407 2489
rect -481 -407 -407 -401
rect 10623 2489 10697 2495
rect 10623 -401 10643 2489
rect 10677 -401 10697 2489
rect 10623 -407 10697 -401
rect -481 -427 10697 -407
rect -481 -461 -401 -427
rect 10617 -461 10697 -427
rect -481 -481 10697 -461
<< nsubdiffcont >>
rect -401 2515 10617 2549
rect -461 -401 -427 2489
rect 10643 -401 10677 2489
rect -401 -461 10617 -427
<< locali >>
rect 102 7501 166 7516
rect 1760 7501 1824 7516
rect 5076 7501 5140 7516
rect 8392 7501 8456 7516
rect 10050 7501 10114 7516
rect -173 7467 -17 7501
rect 102 7467 117 7501
rect 10099 7467 10114 7501
rect 102 7452 166 7467
rect 1760 7452 1824 7467
rect 5076 7452 5140 7467
rect 8392 7452 8456 7467
rect 10050 7452 10114 7467
rect 10739 7501 10803 7516
rect 10739 7467 10754 7501
rect 10788 7467 10803 7501
rect 10739 7452 10803 7467
rect -173 5839 -17 5873
rect 102 5091 166 5106
rect 102 5057 117 5091
rect 151 5057 166 5091
rect 102 5042 166 5057
rect 1760 5091 1824 5106
rect 1760 5057 1775 5091
rect 1809 5057 1824 5091
rect 1760 5042 1824 5057
rect 5076 5091 5140 5106
rect 5076 5057 5091 5091
rect 5125 5057 5140 5091
rect 5076 5042 5140 5057
rect 8392 5091 8456 5106
rect 8392 5057 8407 5091
rect 8441 5057 8456 5091
rect 8392 5042 8456 5057
rect 10050 5091 10114 5106
rect 10050 5057 10065 5091
rect 10099 5057 10114 5091
rect 10050 5042 10114 5057
rect 10739 5453 10803 5468
rect 10739 5419 10754 5453
rect 10788 5419 10803 5453
rect 10739 5404 10803 5419
rect 102 4557 166 4572
rect 5076 4557 5140 4572
rect 10050 4557 10114 4572
rect 102 4523 117 4557
rect 10099 4523 10114 4557
rect 102 4508 166 4523
rect 5076 4508 5140 4523
rect 10050 4508 10114 4523
rect 10421 4406 10485 4421
rect 10421 4288 10436 4406
rect 10470 4288 10485 4406
rect 10421 4273 10485 4288
rect 10945 4406 11009 4421
rect 10945 4288 10960 4406
rect 10994 4288 11009 4406
rect 10945 4273 11009 4288
rect 102 4168 166 4183
rect 1760 4168 1824 4183
rect 5076 4168 5140 4183
rect 8392 4168 8456 4183
rect 10050 4168 10114 4183
rect -203 4134 -17 4168
rect 102 4134 117 4168
rect 10099 4134 10114 4168
rect 102 4119 166 4134
rect 1760 4119 1824 4134
rect 5076 4119 5140 4134
rect 8392 4119 8456 4134
rect 10050 4119 10114 4134
rect 102 3288 166 3303
rect 1760 3288 1824 3303
rect 5076 3288 5140 3303
rect 8392 3288 8456 3303
rect 10050 3288 10114 3303
rect -203 3254 -17 3288
rect 102 3254 117 3288
rect 10099 3254 10114 3288
rect 102 3239 166 3254
rect 1760 3239 1824 3254
rect 5076 3239 5140 3254
rect 8392 3239 8456 3254
rect 10050 3239 10114 3254
rect 1456 2549 1520 2564
rect 5230 2549 5294 2564
rect 8696 2549 8760 2564
rect -461 2515 -401 2549
rect 10617 2515 10677 2549
rect -461 2489 -427 2515
rect 1456 2500 1520 2515
rect 5230 2500 5294 2515
rect 8696 2500 8760 2515
rect 10643 2489 10677 2515
rect 3418 2105 3482 2120
rect 3418 2071 3433 2105
rect 3467 2071 3482 2105
rect 3418 2056 3482 2071
rect 6734 2105 6798 2120
rect 6734 2071 6749 2105
rect 6783 2071 6798 2105
rect 6734 2056 6798 2071
rect 3418 17 3482 32
rect 3418 -17 3433 17
rect 3467 -17 3482 17
rect 3418 -32 3482 -17
rect 6734 16 6798 31
rect 6734 -18 6749 16
rect 6783 -18 6798 16
rect 6734 -33 6798 -18
rect -461 -427 -427 -401
rect 1456 -427 1520 -412
rect 5230 -427 5294 -412
rect 8696 -427 8760 -412
rect 10643 -427 10677 -401
rect -461 -461 -401 -427
rect 10617 -461 10677 -427
rect 1456 -476 1520 -461
rect 5230 -476 5294 -461
rect 8696 -476 8760 -461
<< viali >>
rect 117 7467 10099 7501
rect 10754 7467 10788 7501
rect -17 4598 17 7399
rect 117 5057 151 5091
rect 1775 5057 1809 5091
rect 5091 5057 5125 5091
rect 8407 5057 8441 5091
rect 10065 5057 10099 5091
rect 10199 4646 10233 7447
rect 10754 5419 10788 5453
rect 117 4523 10099 4557
rect 10436 4288 10470 4406
rect 10960 4288 10994 4406
rect 117 4134 10099 4168
rect 117 3254 10099 3288
rect -307 2515 10040 2549
rect -461 -330 -427 2426
rect 3433 2071 3467 2105
rect 6749 2071 6783 2105
rect 3433 -17 3467 17
rect 6749 -18 6783 16
rect 10643 -369 10677 2387
rect 50 -461 10397 -427
<< metal1 >>
rect -32 7510 10252 7516
rect -32 7458 108 7510
rect 160 7501 1766 7510
rect 1818 7501 5082 7510
rect 5134 7501 8398 7510
rect 8450 7501 10056 7510
rect 160 7458 1766 7467
rect 1818 7458 5082 7467
rect 5134 7458 8398 7467
rect 8450 7458 10056 7467
rect 10108 7458 10252 7510
rect -32 7452 10252 7458
rect 10739 7510 10803 7516
rect 10739 7458 10745 7510
rect 10797 7458 10803 7510
rect 10739 7452 10803 7458
rect -32 7399 32 7452
rect -614 7223 -550 7229
rect -614 7171 -608 7223
rect -556 7171 -550 7223
rect -614 7165 -550 7171
rect -356 7223 -292 7229
rect -356 7171 -350 7223
rect -298 7171 -292 7223
rect -356 7165 -292 7171
rect -485 7115 -421 7121
rect -485 7063 -479 7115
rect -427 7063 -421 7115
rect -485 7057 -421 7063
rect -614 6858 -550 6864
rect -614 6806 -608 6858
rect -556 6806 -550 6858
rect -614 6800 -550 6806
rect -356 6858 -292 6864
rect -356 6806 -350 6858
rect -298 6806 -292 6858
rect -356 6800 -292 6806
rect -485 6750 -421 6756
rect -485 6698 -479 6750
rect -427 6698 -421 6750
rect -485 6692 -421 6698
rect -614 6493 -550 6499
rect -614 6441 -608 6493
rect -556 6441 -550 6493
rect -614 6435 -550 6441
rect -356 6481 -292 6487
rect -356 6429 -350 6481
rect -298 6429 -292 6481
rect -356 6423 -292 6429
rect -485 6385 -421 6391
rect -485 6333 -479 6385
rect -427 6333 -421 6385
rect -485 6327 -421 6333
rect -614 6116 -550 6122
rect -614 6064 -608 6116
rect -556 6064 -550 6116
rect -614 6058 -550 6064
rect -356 6116 -292 6122
rect -356 6064 -350 6116
rect -298 6064 -292 6116
rect -356 6058 -292 6064
rect -485 6020 -421 6026
rect -485 5968 -479 6020
rect -427 5968 -421 6020
rect -485 5962 -421 5968
rect -515 5107 -451 5113
rect -515 5055 -509 5107
rect -457 5055 -451 5107
rect -515 5049 -451 5055
rect -644 5020 -580 5026
rect -644 4968 -638 5020
rect -586 4968 -580 5020
rect -644 4962 -580 4968
rect -386 5020 -322 5026
rect -386 4968 -380 5020
rect -328 4968 -322 5020
rect -386 4962 -322 4968
rect -567 4751 -503 4757
rect -567 4699 -561 4751
rect -509 4699 -503 4751
rect -567 4693 -503 4699
rect -386 4664 -322 4670
rect -386 4612 -380 4664
rect -328 4612 -322 4664
rect -386 4606 -322 4612
rect -32 4598 -17 7399
rect 17 4598 32 7399
rect 10188 7447 10252 7452
rect 102 7336 166 7342
rect 102 7284 108 7336
rect 160 7284 166 7336
rect 102 7278 166 7284
rect 1760 7336 1824 7342
rect 1760 7284 1766 7336
rect 1818 7284 1824 7336
rect 1760 7278 1824 7284
rect 3418 7336 3482 7342
rect 3418 7284 3424 7336
rect 3476 7284 3482 7336
rect 3418 7278 3482 7284
rect 5076 7336 5140 7342
rect 5076 7284 5082 7336
rect 5134 7284 5140 7336
rect 5076 7278 5140 7284
rect 6734 7336 6798 7342
rect 6734 7284 6740 7336
rect 6792 7284 6798 7336
rect 6734 7278 6798 7284
rect 8392 7336 8456 7342
rect 8392 7284 8398 7336
rect 8450 7284 8456 7336
rect 8392 7278 8456 7284
rect 10050 7336 10114 7342
rect 10050 7284 10056 7336
rect 10108 7284 10114 7336
rect 10050 7278 10114 7284
rect 111 7227 157 7268
rect 3427 7227 3473 7268
rect 6743 7227 6789 7268
rect 10059 7227 10105 7268
rect 111 7181 167 7227
rect 3417 7181 3483 7227
rect 6733 7181 6799 7227
rect 10049 7181 10105 7227
rect 3427 7093 3473 7181
rect 6743 7093 6789 7181
rect 102 7087 166 7093
rect 102 7035 108 7087
rect 160 7035 166 7087
rect 102 7029 166 7035
rect 1760 7087 1824 7093
rect 1760 7035 1766 7087
rect 1818 7035 1824 7087
rect 1760 7029 1824 7035
rect 3418 7087 3482 7093
rect 3418 7035 3424 7087
rect 3476 7035 3482 7087
rect 3418 7029 3482 7035
rect 5076 7087 5140 7093
rect 5076 7035 5082 7087
rect 5134 7035 5140 7087
rect 5076 7029 5140 7035
rect 6734 7087 6798 7093
rect 6734 7035 6740 7087
rect 6792 7035 6798 7087
rect 6734 7029 6798 7035
rect 8392 7087 8456 7093
rect 8392 7035 8398 7087
rect 8450 7035 8456 7087
rect 8392 7029 8456 7035
rect 10050 7087 10114 7093
rect 10050 7035 10056 7087
rect 10108 7035 10114 7087
rect 10050 7029 10114 7035
rect 111 6978 157 7019
rect 3427 6978 3473 7029
rect 6743 6978 6789 7029
rect 10059 6978 10105 7019
rect 111 6932 167 6978
rect 3417 6932 3483 6978
rect 6733 6932 6799 6978
rect 10049 6932 10105 6978
rect 3427 6844 3473 6932
rect 6743 6844 6789 6932
rect 102 6838 166 6844
rect 102 6786 108 6838
rect 160 6786 166 6838
rect 102 6780 166 6786
rect 1760 6838 1824 6844
rect 1760 6786 1766 6838
rect 1818 6786 1824 6838
rect 1760 6780 1824 6786
rect 3418 6838 3482 6844
rect 3418 6786 3424 6838
rect 3476 6786 3482 6838
rect 3418 6780 3482 6786
rect 5076 6838 5140 6844
rect 5076 6786 5082 6838
rect 5134 6786 5140 6838
rect 5076 6780 5140 6786
rect 6734 6838 6798 6844
rect 6734 6786 6740 6838
rect 6792 6786 6798 6838
rect 6734 6780 6798 6786
rect 8392 6838 8456 6844
rect 8392 6786 8398 6838
rect 8450 6786 8456 6838
rect 8392 6780 8456 6786
rect 10050 6838 10114 6844
rect 10050 6786 10056 6838
rect 10108 6786 10114 6838
rect 10050 6780 10114 6786
rect 111 6729 157 6770
rect 3427 6729 3473 6780
rect 6743 6729 6789 6780
rect 10059 6729 10105 6770
rect 111 6683 167 6729
rect 3417 6683 3483 6729
rect 6733 6683 6799 6729
rect 10049 6683 10105 6729
rect 3427 6595 3473 6683
rect 6743 6595 6789 6683
rect 102 6589 166 6595
rect 102 6537 108 6589
rect 160 6537 166 6589
rect 102 6531 166 6537
rect 1760 6589 1824 6595
rect 1760 6537 1766 6589
rect 1818 6537 1824 6589
rect 1760 6531 1824 6537
rect 3418 6589 3482 6595
rect 3418 6537 3424 6589
rect 3476 6537 3482 6589
rect 3418 6531 3482 6537
rect 5076 6589 5140 6595
rect 5076 6537 5082 6589
rect 5134 6537 5140 6589
rect 5076 6531 5140 6537
rect 6734 6589 6798 6595
rect 6734 6537 6740 6589
rect 6792 6537 6798 6589
rect 6734 6531 6798 6537
rect 8392 6589 8456 6595
rect 8392 6537 8398 6589
rect 8450 6537 8456 6589
rect 8392 6531 8456 6537
rect 10050 6589 10114 6595
rect 10050 6537 10056 6589
rect 10108 6537 10114 6589
rect 10050 6531 10114 6537
rect 111 6480 157 6521
rect 3427 6480 3473 6531
rect 6743 6480 6789 6531
rect 10059 6480 10105 6521
rect 111 6434 167 6480
rect 3417 6434 3483 6480
rect 6733 6434 6799 6480
rect 10049 6434 10105 6480
rect 102 6340 166 6346
rect 102 6288 108 6340
rect 160 6288 166 6340
rect 102 6282 166 6288
rect 1760 6340 1824 6346
rect 1760 6288 1766 6340
rect 1818 6288 1824 6340
rect 1760 6282 1824 6288
rect 3418 6340 3482 6346
rect 3418 6288 3424 6340
rect 3476 6288 3482 6340
rect 3418 6282 3482 6288
rect 5076 6340 5140 6346
rect 5076 6288 5082 6340
rect 5134 6288 5140 6340
rect 5076 6282 5140 6288
rect 6734 6340 6798 6346
rect 6734 6288 6740 6340
rect 6792 6288 6798 6340
rect 6734 6282 6798 6288
rect 8392 6340 8456 6346
rect 8392 6288 8398 6340
rect 8450 6288 8456 6340
rect 8392 6282 8456 6288
rect 10050 6340 10114 6346
rect 10050 6288 10056 6340
rect 10108 6288 10114 6340
rect 10050 6282 10114 6288
rect 111 6231 157 6272
rect 4300 6234 4364 6240
rect 111 6185 167 6231
rect 3417 6185 3483 6231
rect 4300 6182 4306 6234
rect 4358 6182 4364 6234
rect 4300 6176 4364 6182
rect 5956 6234 6020 6240
rect 5956 6182 5962 6234
rect 6014 6182 6020 6234
rect 10059 6231 10105 6272
rect 6733 6185 6799 6231
rect 10049 6185 10105 6231
rect 5956 6176 6020 6182
rect 102 6091 166 6097
rect 102 6039 108 6091
rect 160 6039 166 6091
rect 102 6033 166 6039
rect 1760 6091 1824 6097
rect 1760 6039 1766 6091
rect 1818 6039 1824 6091
rect 1760 6033 1824 6039
rect 3418 6091 3482 6097
rect 3418 6039 3424 6091
rect 3476 6039 3482 6091
rect 3418 6033 3482 6039
rect 5076 6091 5140 6097
rect 5076 6039 5082 6091
rect 5134 6039 5140 6091
rect 5076 6033 5140 6039
rect 6734 6091 6798 6097
rect 6734 6039 6740 6091
rect 6792 6039 6798 6091
rect 6734 6033 6798 6039
rect 8392 6091 8456 6097
rect 8392 6039 8398 6091
rect 8450 6039 8456 6091
rect 8392 6033 8456 6039
rect 10050 6091 10114 6097
rect 10050 6039 10056 6091
rect 10108 6039 10114 6091
rect 10050 6033 10114 6039
rect 111 5982 157 6023
rect 4300 5985 4364 5991
rect 111 5936 167 5982
rect 3417 5936 3483 5982
rect 4300 5933 4306 5985
rect 4358 5933 4364 5985
rect 4300 5927 4364 5933
rect 5956 5985 6020 5991
rect 5956 5933 5962 5985
rect 6014 5933 6020 5985
rect 10059 5982 10105 6023
rect 6733 5936 6799 5982
rect 10049 5936 10105 5982
rect 5956 5927 6020 5933
rect 102 5842 166 5848
rect 102 5790 108 5842
rect 160 5790 166 5842
rect 102 5784 166 5790
rect 1760 5842 1824 5848
rect 1760 5790 1766 5842
rect 1818 5790 1824 5842
rect 1760 5784 1824 5790
rect 3418 5842 3482 5848
rect 3418 5790 3424 5842
rect 3476 5790 3482 5842
rect 3418 5784 3482 5790
rect 5076 5842 5140 5848
rect 5076 5790 5082 5842
rect 5134 5790 5140 5842
rect 5076 5784 5140 5790
rect 6734 5842 6798 5848
rect 6734 5790 6740 5842
rect 6792 5790 6798 5842
rect 6734 5784 6798 5790
rect 8392 5842 8456 5848
rect 8392 5790 8398 5842
rect 8450 5790 8456 5842
rect 8392 5784 8456 5790
rect 10050 5842 10114 5848
rect 10050 5790 10056 5842
rect 10108 5790 10114 5842
rect 10050 5784 10114 5790
rect 111 5733 157 5774
rect 4300 5736 4364 5742
rect 111 5687 167 5733
rect 3417 5687 3483 5733
rect 4300 5684 4306 5736
rect 4358 5684 4364 5736
rect 4300 5678 4364 5684
rect 5956 5736 6020 5742
rect 5956 5684 5962 5736
rect 6014 5684 6020 5736
rect 10059 5733 10105 5774
rect 6733 5687 6799 5733
rect 10049 5687 10105 5733
rect 5956 5678 6020 5684
rect 102 5593 166 5599
rect 102 5541 108 5593
rect 160 5541 166 5593
rect 102 5535 166 5541
rect 1760 5593 1824 5599
rect 1760 5541 1766 5593
rect 1818 5541 1824 5593
rect 1760 5535 1824 5541
rect 3418 5593 3482 5599
rect 3418 5541 3424 5593
rect 3476 5541 3482 5593
rect 3418 5535 3482 5541
rect 5076 5593 5140 5599
rect 5076 5541 5082 5593
rect 5134 5541 5140 5593
rect 5076 5535 5140 5541
rect 6734 5593 6798 5599
rect 6734 5541 6740 5593
rect 6792 5541 6798 5593
rect 6734 5535 6798 5541
rect 8392 5593 8456 5599
rect 8392 5541 8398 5593
rect 8450 5541 8456 5593
rect 8392 5535 8456 5541
rect 10050 5593 10114 5599
rect 10050 5541 10056 5593
rect 10108 5541 10114 5593
rect 10050 5535 10114 5541
rect 111 5484 157 5525
rect 4300 5487 4364 5493
rect 111 5438 167 5484
rect 3417 5438 3483 5484
rect 4300 5435 4306 5487
rect 4358 5435 4364 5487
rect 4300 5429 4364 5435
rect 5956 5487 6020 5493
rect 5956 5435 5962 5487
rect 6014 5435 6020 5487
rect 10059 5484 10105 5525
rect 6733 5438 6799 5484
rect 10049 5438 10105 5484
rect 5956 5429 6020 5435
rect 102 5344 166 5350
rect 102 5292 108 5344
rect 160 5292 166 5344
rect 102 5286 166 5292
rect 1760 5344 1824 5350
rect 1760 5292 1766 5344
rect 1818 5292 1824 5344
rect 1760 5286 1824 5292
rect 3418 5344 3482 5350
rect 3418 5292 3424 5344
rect 3476 5292 3482 5344
rect 3418 5286 3482 5292
rect 5076 5344 5140 5350
rect 5076 5292 5082 5344
rect 5134 5292 5140 5344
rect 5076 5286 5140 5292
rect 6734 5344 6798 5350
rect 6734 5292 6740 5344
rect 6792 5292 6798 5344
rect 6734 5286 6798 5292
rect 8392 5344 8456 5350
rect 8392 5292 8398 5344
rect 8450 5292 8456 5344
rect 8392 5286 8456 5292
rect 10050 5344 10114 5350
rect 10050 5292 10056 5344
rect 10108 5292 10114 5344
rect 10050 5286 10114 5292
rect 111 5235 157 5276
rect 4300 5238 4364 5244
rect 111 5189 167 5235
rect 3417 5189 3483 5235
rect 4300 5186 4306 5238
rect 4358 5186 4364 5238
rect 4300 5180 4364 5186
rect 5956 5238 6020 5244
rect 5956 5186 5962 5238
rect 6014 5186 6020 5238
rect 10059 5235 10105 5276
rect 6733 5189 6799 5235
rect 10049 5189 10105 5235
rect 5956 5180 6020 5186
rect 102 5100 166 5106
rect 102 5048 108 5100
rect 160 5048 166 5100
rect 102 5042 166 5048
rect 1760 5100 1824 5106
rect 1760 5048 1766 5100
rect 1818 5048 1824 5100
rect 1760 5042 1824 5048
rect 5076 5100 5140 5106
rect 5076 5048 5082 5100
rect 5134 5048 5140 5100
rect 5076 5042 5140 5048
rect 8392 5100 8456 5106
rect 8392 5048 8398 5100
rect 8450 5048 8456 5100
rect 8392 5042 8456 5048
rect 10050 5100 10114 5106
rect 10050 5048 10056 5100
rect 10108 5048 10114 5100
rect 10050 5042 10114 5048
rect 102 4937 166 4943
rect 102 4885 108 4937
rect 160 4885 166 4937
rect 102 4879 166 4885
rect 1760 4937 1824 4943
rect 1760 4885 1766 4937
rect 1818 4885 1824 4937
rect 1760 4879 1824 4885
rect 5076 4937 5140 4943
rect 5076 4885 5082 4937
rect 5134 4885 5140 4937
rect 5076 4879 5140 4885
rect 8392 4937 8456 4943
rect 8392 4885 8398 4937
rect 8450 4885 8456 4937
rect 8392 4879 8456 4885
rect 10050 4937 10114 4943
rect 10050 4885 10056 4937
rect 10108 4885 10114 4937
rect 10050 4879 10114 4885
rect 3418 4807 3482 4813
rect 3418 4755 3424 4807
rect 3476 4755 3482 4807
rect 3418 4749 3482 4755
rect 6734 4807 6798 4813
rect 6734 4755 6740 4807
rect 6792 4755 6798 4807
rect 6734 4749 6798 4755
rect 111 4702 157 4743
rect 4300 4705 4364 4711
rect 111 4656 167 4702
rect 3417 4656 3483 4702
rect 4300 4653 4306 4705
rect 4358 4653 4364 4705
rect 4300 4647 4364 4653
rect 5956 4705 6020 4711
rect 5956 4653 5962 4705
rect 6014 4653 6020 4705
rect 10059 4702 10105 4743
rect 6733 4656 6799 4702
rect 10049 4656 10105 4702
rect 5956 4647 6020 4653
rect -32 4572 32 4598
rect 10188 4646 10199 7447
rect 10233 4646 10252 7447
rect 10739 7376 10803 7382
rect 10739 7324 10745 7376
rect 10797 7324 10803 7376
rect 10739 7318 10803 7324
rect 10522 6071 10568 7205
rect 10609 7198 10673 7204
rect 10609 7146 10615 7198
rect 10667 7146 10673 7198
rect 10609 7140 10673 7146
rect 10739 7020 10803 7026
rect 10739 6968 10745 7020
rect 10797 6968 10803 7020
rect 10739 6962 10803 6968
rect 10609 6842 10673 6848
rect 10609 6790 10615 6842
rect 10667 6790 10673 6842
rect 10609 6784 10673 6790
rect 10739 6664 10803 6670
rect 10739 6612 10745 6664
rect 10797 6612 10803 6664
rect 10739 6606 10803 6612
rect 10609 6486 10673 6492
rect 10609 6434 10615 6486
rect 10667 6434 10673 6486
rect 10609 6428 10673 6434
rect 10739 6308 10803 6314
rect 10739 6256 10745 6308
rect 10797 6256 10803 6308
rect 10739 6250 10803 6256
rect 10609 6130 10673 6136
rect 10609 6078 10615 6130
rect 10667 6078 10673 6130
rect 10609 6072 10673 6078
rect 10506 6007 10570 6013
rect 10506 5955 10512 6007
rect 10564 5955 10570 6007
rect 10506 5949 10570 5955
rect 10739 5952 10803 5958
rect 10739 5900 10745 5952
rect 10797 5900 10803 5952
rect 10739 5894 10803 5900
rect 10522 5715 10568 5781
rect 10609 5774 10673 5780
rect 10609 5722 10615 5774
rect 10667 5722 10673 5774
rect 10609 5716 10673 5722
rect 10508 5661 10572 5667
rect 10508 5609 10514 5661
rect 10566 5609 10572 5661
rect 10508 5603 10572 5609
rect 10739 5596 10803 5602
rect 10739 5544 10745 5596
rect 10797 5544 10803 5596
rect 10739 5538 10803 5544
rect 10739 5462 10803 5468
rect 10739 5410 10745 5462
rect 10797 5410 10803 5462
rect 10739 5404 10803 5410
rect 10774 5096 10838 5102
rect 10774 5044 10780 5096
rect 10832 5044 10838 5096
rect 10774 5038 10838 5044
rect 10188 4572 10252 4646
rect -32 4566 10252 4572
rect -644 4528 -580 4534
rect -644 4476 -638 4528
rect -586 4476 -580 4528
rect -32 4514 108 4566
rect 160 4557 1766 4566
rect 1818 4557 5082 4566
rect 5134 4557 10056 4566
rect 160 4514 1766 4523
rect 1818 4514 5082 4523
rect 5134 4514 10056 4523
rect 10108 4514 10252 4566
rect -32 4508 10252 4514
rect -644 4470 -580 4476
rect 10421 4415 10485 4421
rect -515 4395 -451 4401
rect -515 4343 -509 4395
rect -457 4343 -451 4395
rect -515 4337 -451 4343
rect 10421 4279 10427 4415
rect 10479 4279 10485 4415
rect 10421 4273 10485 4279
rect -386 4184 -322 4190
rect -644 4172 -580 4178
rect -644 4120 -638 4172
rect -586 4120 -580 4172
rect -386 4132 -380 4184
rect -328 4132 -322 4184
rect -386 4126 -322 4132
rect -32 4177 10248 4183
rect -644 4114 -580 4120
rect -32 4125 108 4177
rect 160 4168 1766 4177
rect 1818 4168 5082 4177
rect 5134 4168 8398 4177
rect 8450 4168 10056 4177
rect 160 4125 1766 4134
rect 1818 4125 5082 4134
rect 5134 4125 8398 4134
rect 8450 4125 10056 4134
rect 10108 4125 10248 4177
rect -32 4119 10248 4125
rect -515 4039 -451 4045
rect -515 3987 -509 4039
rect -457 3987 -451 4039
rect -515 3981 -451 3987
rect -386 3952 -322 3958
rect -386 3900 -380 3952
rect -328 3900 -322 3952
rect -386 3894 -322 3900
rect -644 3816 -580 3822
rect -644 3764 -638 3816
rect -586 3764 -580 3816
rect -644 3758 -580 3764
rect -515 3683 -451 3689
rect -515 3631 -509 3683
rect -457 3631 -451 3683
rect -515 3625 -451 3631
rect -386 3596 -322 3602
rect -386 3544 -380 3596
rect -327 3544 -322 3596
rect -386 3538 -322 3544
rect -644 3460 -580 3466
rect -644 3408 -638 3460
rect -586 3408 -580 3460
rect -644 3402 -580 3408
rect -32 3303 32 4119
rect 108 3990 167 4036
rect 3417 3990 3483 4036
rect 5075 3990 5141 4036
rect 6733 3990 6799 4036
rect 10049 3990 10108 4036
rect 108 3952 160 3990
rect 3427 3952 3473 3990
rect 10056 3952 10108 3990
rect 102 3946 166 3952
rect 102 3894 108 3946
rect 160 3894 166 3946
rect 102 3888 166 3894
rect 1760 3946 1824 3952
rect 1760 3894 1766 3946
rect 1818 3894 1824 3946
rect 1760 3888 1824 3894
rect 3418 3946 3482 3952
rect 3418 3894 3424 3946
rect 3476 3894 3482 3946
rect 3418 3888 3482 3894
rect 5076 3946 5140 3952
rect 5076 3894 5082 3946
rect 5134 3894 5140 3946
rect 5076 3888 5140 3894
rect 6734 3947 6798 3952
rect 6734 3894 6740 3947
rect 6792 3894 6798 3947
rect 6734 3888 6798 3894
rect 8392 3946 8456 3952
rect 8392 3894 8398 3946
rect 8450 3894 8456 3946
rect 8392 3888 8456 3894
rect 10050 3946 10114 3952
rect 10050 3894 10056 3946
rect 10108 3894 10114 3946
rect 10050 3888 10114 3894
rect 108 3634 167 3680
rect 3417 3634 3483 3680
rect 5075 3634 5141 3680
rect 6733 3634 6799 3680
rect 10049 3634 10108 3680
rect 108 3596 160 3634
rect 3427 3596 3473 3634
rect 10056 3596 10108 3634
rect 102 3590 166 3596
rect 102 3538 108 3590
rect 160 3538 166 3590
rect 102 3532 166 3538
rect 1760 3590 1824 3596
rect 1760 3538 1766 3590
rect 1818 3538 1824 3590
rect 1760 3532 1824 3538
rect 3418 3590 3482 3596
rect 3418 3538 3424 3590
rect 3476 3538 3482 3590
rect 3418 3532 3482 3538
rect 5076 3590 5140 3596
rect 5076 3538 5082 3590
rect 5134 3538 5140 3590
rect 5076 3532 5140 3538
rect 8392 3590 8456 3596
rect 8392 3538 8398 3590
rect 8450 3538 8456 3590
rect 8392 3532 8456 3538
rect 10050 3590 10114 3596
rect 10050 3538 10056 3590
rect 10108 3538 10114 3590
rect 10050 3532 10114 3538
rect 6734 3466 6798 3472
rect 6734 3414 6740 3466
rect 6792 3414 6798 3466
rect 6734 3408 6798 3414
rect 10184 3303 10248 4119
rect 10560 3791 10606 4925
rect 10643 4919 10707 4925
rect 10643 4867 10649 4919
rect 10701 4867 10707 4919
rect 10643 4861 10707 4867
rect 10774 4740 10838 4746
rect 10774 4688 10780 4740
rect 10832 4688 10838 4740
rect 10774 4682 10838 4688
rect 10643 4563 10707 4569
rect 10643 4511 10649 4563
rect 10701 4511 10707 4563
rect 10643 4505 10707 4511
rect 10945 4415 11009 4421
rect 10774 4384 10838 4390
rect 10774 4332 10780 4384
rect 10832 4332 10838 4384
rect 10774 4326 10838 4332
rect 10945 4279 10951 4415
rect 11003 4279 11009 4415
rect 10945 4273 11009 4279
rect 10643 4207 10707 4213
rect 10643 4155 10649 4207
rect 10701 4155 10707 4207
rect 10643 4149 10707 4155
rect 10774 4028 10838 4034
rect 10774 3976 10780 4028
rect 10832 3976 10838 4028
rect 10774 3970 10838 3976
rect 10643 3851 10707 3857
rect 10643 3799 10649 3851
rect 10701 3799 10707 3851
rect 10643 3793 10707 3799
rect 10539 3728 10603 3734
rect 10539 3676 10545 3728
rect 10597 3676 10603 3728
rect 10539 3670 10603 3676
rect 10774 3672 10838 3678
rect 10774 3620 10780 3672
rect 10832 3620 10838 3672
rect 10774 3614 10838 3620
rect 10545 3608 10609 3614
rect 10545 3556 10551 3608
rect 10603 3556 10609 3608
rect 10545 3550 10609 3556
rect 10560 3435 10606 3501
rect 10645 3494 10709 3500
rect 10645 3442 10651 3494
rect 10703 3442 10709 3494
rect 10645 3436 10709 3442
rect -32 3297 10248 3303
rect -32 3245 108 3297
rect 160 3288 1766 3297
rect 1818 3288 5082 3297
rect 5134 3288 8398 3297
rect 8450 3288 10056 3297
rect 160 3245 1766 3254
rect 1818 3245 5082 3254
rect 5134 3245 8398 3254
rect 8450 3245 10056 3254
rect 10108 3245 10248 3297
rect 10774 3316 10838 3322
rect 10774 3264 10780 3316
rect 10832 3264 10838 3316
rect 10774 3258 10838 3264
rect -32 3239 10248 3245
rect -476 2558 10692 2564
rect -476 2549 1462 2558
rect 1514 2549 5236 2558
rect 5288 2549 8702 2558
rect 8754 2549 10692 2558
rect -476 2515 -307 2549
rect 10040 2515 10692 2549
rect -476 2506 1462 2515
rect 1514 2506 5236 2515
rect 5288 2506 8702 2515
rect 8754 2506 10692 2515
rect -476 2500 10692 2506
rect -476 2426 -412 2500
rect -476 -330 -461 2426
rect -427 -330 -412 2426
rect 10628 2387 10692 2500
rect 3418 2114 3482 2120
rect 3418 2062 3424 2114
rect 3476 2062 3482 2114
rect 3418 2056 3482 2062
rect 6734 2114 6798 2120
rect 6734 2062 6740 2114
rect 6792 2062 6798 2114
rect 6734 2056 6798 2062
rect 3138 1976 3202 1982
rect 3138 1924 3144 1976
rect 3196 1924 3202 1976
rect 3138 1918 3202 1924
rect 4725 1976 4789 1982
rect 4725 1924 4731 1976
rect 4783 1924 4789 1976
rect 6957 1976 7021 1982
rect 5075 1927 5141 1973
rect 4725 1918 4789 1924
rect 6957 1924 6963 1976
rect 7015 1924 7021 1976
rect 6957 1918 7021 1924
rect 102 1827 108 1879
rect 160 1827 166 1879
rect 1760 1827 1766 1879
rect 1818 1827 1824 1879
rect 3418 1827 3424 1879
rect 3476 1827 3482 1879
rect 5076 1827 5082 1879
rect 5134 1827 5140 1879
rect 6734 1827 6740 1879
rect 6792 1827 6798 1879
rect 8392 1827 8398 1879
rect 8450 1827 8456 1879
rect 10050 1827 10056 1879
rect 10108 1827 10114 1879
rect 3138 1736 3202 1742
rect 3138 1684 3144 1736
rect 3196 1684 3202 1736
rect 3138 1678 3202 1684
rect 4725 1736 4789 1742
rect 4725 1684 4731 1736
rect 4783 1684 4789 1736
rect 6957 1736 7021 1742
rect 5075 1687 5141 1733
rect 4725 1678 4789 1684
rect 6957 1684 6963 1736
rect 7015 1684 7021 1736
rect 6957 1678 7021 1684
rect 102 1587 108 1639
rect 160 1587 166 1639
rect 1760 1587 1766 1639
rect 1818 1587 1824 1639
rect 3418 1587 3424 1639
rect 3476 1587 3482 1639
rect 5076 1587 5082 1639
rect 5134 1587 5140 1639
rect 6734 1587 6740 1639
rect 6792 1587 6798 1639
rect 8392 1587 8398 1639
rect 8450 1587 8456 1639
rect 10050 1587 10056 1639
rect 10108 1587 10114 1639
rect 3138 1496 3202 1502
rect 3138 1444 3144 1496
rect 3196 1444 3202 1496
rect 3138 1438 3202 1444
rect 4725 1496 4789 1502
rect 4725 1444 4731 1496
rect 4783 1444 4789 1496
rect 6957 1496 7021 1502
rect 5075 1447 5141 1493
rect 4725 1438 4789 1444
rect 6957 1444 6963 1496
rect 7015 1444 7021 1496
rect 6957 1438 7021 1444
rect 102 1347 108 1399
rect 160 1347 166 1399
rect 1760 1347 1766 1399
rect 1818 1347 1824 1399
rect 3418 1347 3424 1399
rect 3476 1347 3482 1399
rect 5076 1347 5082 1399
rect 5134 1347 5140 1399
rect 6734 1347 6740 1399
rect 6792 1347 6798 1399
rect 8392 1347 8398 1399
rect 8450 1347 8456 1399
rect 10050 1347 10056 1399
rect 10108 1347 10114 1399
rect 3138 1256 3202 1262
rect 3138 1204 3144 1256
rect 3196 1204 3202 1256
rect 3138 1198 3202 1204
rect 4725 1256 4789 1262
rect 4725 1204 4731 1256
rect 4783 1204 4789 1256
rect 6957 1256 7021 1262
rect 5075 1207 5141 1253
rect 4725 1198 4789 1204
rect 6957 1204 6963 1256
rect 7015 1204 7021 1256
rect 6957 1198 7021 1204
rect 102 1107 108 1159
rect 160 1107 166 1159
rect 1760 1107 1766 1159
rect 1818 1107 1824 1159
rect 3418 1107 3424 1159
rect 3476 1107 3482 1159
rect 5076 1107 5082 1159
rect 5134 1107 5140 1159
rect 6734 1107 6740 1159
rect 6792 1107 6798 1159
rect 8392 1107 8398 1159
rect 8450 1107 8456 1159
rect 10050 1107 10056 1159
rect 10108 1107 10114 1159
rect 3138 1016 3202 1022
rect 3138 964 3144 1016
rect 3196 964 3202 1016
rect 3138 958 3202 964
rect 4725 1016 4789 1022
rect 4725 964 4731 1016
rect 4783 964 4789 1016
rect 6957 1016 7021 1022
rect 5075 967 5141 1013
rect 4725 958 4789 964
rect 6957 964 6963 1016
rect 7015 964 7021 1016
rect 6957 958 7021 964
rect 102 867 108 919
rect 160 867 166 919
rect 1760 867 1766 919
rect 1818 867 1824 919
rect 3418 867 3424 919
rect 3476 867 3482 919
rect 5076 867 5082 919
rect 5134 867 5140 919
rect 6734 867 6740 919
rect 6792 867 6798 919
rect 8392 867 8398 919
rect 8450 867 8456 919
rect 10050 867 10056 919
rect 10108 867 10114 919
rect 3138 776 3202 782
rect 3138 724 3144 776
rect 3196 724 3202 776
rect 3138 718 3202 724
rect 4725 776 4789 782
rect 4725 724 4731 776
rect 4783 724 4789 776
rect 6957 776 7021 782
rect 5075 727 5141 773
rect 4725 718 4789 724
rect 6957 724 6963 776
rect 7015 724 7021 776
rect 6957 718 7021 724
rect 102 627 108 679
rect 160 627 166 679
rect 1760 627 1766 679
rect 1818 627 1824 679
rect 3418 627 3424 679
rect 3476 627 3482 679
rect 5076 627 5082 679
rect 5134 627 5140 679
rect 6734 627 6740 679
rect 6792 627 6798 679
rect 8392 627 8398 679
rect 8450 627 8456 679
rect 10050 627 10056 679
rect 10108 627 10114 679
rect 3138 536 3202 542
rect 3138 484 3144 536
rect 3196 484 3202 536
rect 3138 478 3202 484
rect 4725 536 4789 542
rect 4725 484 4731 536
rect 4783 484 4789 536
rect 6957 536 7021 542
rect 5075 487 5141 533
rect 4725 478 4789 484
rect 6957 484 6963 536
rect 7015 484 7021 536
rect 6957 478 7021 484
rect 102 387 108 439
rect 160 387 166 439
rect 1760 387 1766 439
rect 1818 387 1824 439
rect 3418 387 3424 439
rect 3476 387 3482 439
rect 5076 387 5082 439
rect 5134 387 5140 439
rect 6734 387 6740 439
rect 6792 387 6798 439
rect 8392 387 8398 439
rect 8450 387 8456 439
rect 10050 387 10056 439
rect 10108 387 10114 439
rect 3138 296 3202 302
rect 3138 244 3144 296
rect 3196 244 3202 296
rect 3138 238 3202 244
rect 4725 296 4789 302
rect 4725 244 4731 296
rect 4783 244 4789 296
rect 6957 296 7021 302
rect 5075 247 5141 293
rect 4725 238 4789 244
rect 6957 244 6963 296
rect 7015 244 7021 296
rect 6957 238 7021 244
rect 102 147 108 199
rect 160 147 166 199
rect 1760 147 1766 199
rect 1818 147 1824 199
rect 3418 147 3424 199
rect 3476 147 3482 199
rect 5076 147 5082 199
rect 5134 147 5140 199
rect 6734 147 6740 199
rect 6792 147 6798 199
rect 8392 147 8398 199
rect 8450 147 8456 199
rect 10050 147 10056 199
rect 10108 147 10114 199
rect 3418 26 3482 32
rect 3418 -26 3424 26
rect 3476 -26 3482 26
rect 3418 -32 3482 -26
rect 6734 25 6798 31
rect 6734 -27 6740 25
rect 6792 -27 6798 25
rect 6734 -33 6798 -27
rect -476 -412 -412 -330
rect 10628 -369 10643 2387
rect 10677 -369 10692 2387
rect 10628 -412 10692 -369
rect -476 -418 10692 -412
rect -476 -427 1462 -418
rect 1514 -427 5236 -418
rect 5288 -427 8702 -418
rect 8754 -427 10692 -418
rect -476 -461 50 -427
rect 10397 -461 10692 -427
rect -476 -470 1462 -461
rect 1514 -470 5236 -461
rect 5288 -470 8702 -461
rect 8754 -470 10692 -461
rect -476 -476 10692 -470
<< via1 >>
rect 108 7501 160 7510
rect 1766 7501 1818 7510
rect 5082 7501 5134 7510
rect 8398 7501 8450 7510
rect 10056 7501 10108 7510
rect 108 7467 117 7501
rect 117 7467 160 7501
rect 1766 7467 1818 7501
rect 5082 7467 5134 7501
rect 8398 7467 8450 7501
rect 10056 7467 10099 7501
rect 10099 7467 10108 7501
rect 108 7458 160 7467
rect 1766 7458 1818 7467
rect 5082 7458 5134 7467
rect 8398 7458 8450 7467
rect 10056 7458 10108 7467
rect 10745 7501 10797 7510
rect 10745 7467 10754 7501
rect 10754 7467 10788 7501
rect 10788 7467 10797 7501
rect 10745 7458 10797 7467
rect -608 7171 -556 7223
rect -350 7171 -298 7223
rect -479 7063 -427 7115
rect -608 6806 -556 6858
rect -350 6806 -298 6858
rect -479 6698 -427 6750
rect -608 6441 -556 6493
rect -350 6429 -298 6481
rect -479 6333 -427 6385
rect -608 6064 -556 6116
rect -350 6064 -298 6116
rect -479 5968 -427 6020
rect -509 5055 -457 5107
rect -638 4968 -586 5020
rect -380 4968 -328 5020
rect -561 4699 -509 4751
rect -380 4612 -328 4664
rect 108 7284 160 7336
rect 1766 7284 1818 7336
rect 3424 7284 3476 7336
rect 5082 7284 5134 7336
rect 6740 7284 6792 7336
rect 8398 7284 8450 7336
rect 10056 7284 10108 7336
rect 108 7035 160 7087
rect 1766 7035 1818 7087
rect 3424 7035 3476 7087
rect 5082 7035 5134 7087
rect 6740 7035 6792 7087
rect 8398 7035 8450 7087
rect 10056 7035 10108 7087
rect 108 6786 160 6838
rect 1766 6786 1818 6838
rect 3424 6786 3476 6838
rect 5082 6786 5134 6838
rect 6740 6786 6792 6838
rect 8398 6786 8450 6838
rect 10056 6786 10108 6838
rect 108 6537 160 6589
rect 1766 6537 1818 6589
rect 3424 6537 3476 6589
rect 5082 6537 5134 6589
rect 6740 6537 6792 6589
rect 8398 6537 8450 6589
rect 10056 6537 10108 6589
rect 108 6288 160 6340
rect 1766 6288 1818 6340
rect 3424 6288 3476 6340
rect 5082 6288 5134 6340
rect 6740 6288 6792 6340
rect 8398 6288 8450 6340
rect 10056 6288 10108 6340
rect 4306 6182 4358 6234
rect 5962 6182 6014 6234
rect 108 6039 160 6091
rect 1766 6039 1818 6091
rect 3424 6039 3476 6091
rect 5082 6039 5134 6091
rect 6740 6039 6792 6091
rect 8398 6039 8450 6091
rect 10056 6039 10108 6091
rect 4306 5933 4358 5985
rect 5962 5933 6014 5985
rect 108 5790 160 5842
rect 1766 5790 1818 5842
rect 3424 5790 3476 5842
rect 5082 5790 5134 5842
rect 6740 5790 6792 5842
rect 8398 5790 8450 5842
rect 10056 5790 10108 5842
rect 4306 5684 4358 5736
rect 5962 5684 6014 5736
rect 108 5541 160 5593
rect 1766 5541 1818 5593
rect 3424 5541 3476 5593
rect 5082 5541 5134 5593
rect 6740 5541 6792 5593
rect 8398 5541 8450 5593
rect 10056 5541 10108 5593
rect 4306 5435 4358 5487
rect 5962 5435 6014 5487
rect 108 5292 160 5344
rect 1766 5292 1818 5344
rect 3424 5292 3476 5344
rect 5082 5292 5134 5344
rect 6740 5292 6792 5344
rect 8398 5292 8450 5344
rect 10056 5292 10108 5344
rect 4306 5186 4358 5238
rect 5962 5186 6014 5238
rect 108 5091 160 5100
rect 108 5057 117 5091
rect 117 5057 151 5091
rect 151 5057 160 5091
rect 108 5048 160 5057
rect 1766 5091 1818 5100
rect 1766 5057 1775 5091
rect 1775 5057 1809 5091
rect 1809 5057 1818 5091
rect 1766 5048 1818 5057
rect 5082 5091 5134 5100
rect 5082 5057 5091 5091
rect 5091 5057 5125 5091
rect 5125 5057 5134 5091
rect 5082 5048 5134 5057
rect 8398 5091 8450 5100
rect 8398 5057 8407 5091
rect 8407 5057 8441 5091
rect 8441 5057 8450 5091
rect 8398 5048 8450 5057
rect 10056 5091 10108 5100
rect 10056 5057 10065 5091
rect 10065 5057 10099 5091
rect 10099 5057 10108 5091
rect 10056 5048 10108 5057
rect 108 4885 160 4937
rect 1766 4885 1818 4937
rect 5082 4885 5134 4937
rect 8398 4885 8450 4937
rect 10056 4885 10108 4937
rect 3424 4755 3476 4807
rect 6740 4755 6792 4807
rect 4306 4653 4358 4705
rect 5962 4653 6014 4705
rect 10745 7324 10797 7376
rect 10615 7146 10667 7198
rect 10745 6968 10797 7020
rect 10615 6790 10667 6842
rect 10745 6612 10797 6664
rect 10615 6434 10667 6486
rect 10745 6256 10797 6308
rect 10615 6078 10667 6130
rect 10512 5955 10564 6007
rect 10745 5900 10797 5952
rect 10615 5722 10667 5774
rect 10514 5609 10566 5661
rect 10745 5544 10797 5596
rect 10745 5453 10797 5462
rect 10745 5419 10754 5453
rect 10754 5419 10788 5453
rect 10788 5419 10797 5453
rect 10745 5410 10797 5419
rect 10780 5044 10832 5096
rect -638 4476 -586 4528
rect 108 4557 160 4566
rect 1766 4557 1818 4566
rect 5082 4557 5134 4566
rect 10056 4557 10108 4566
rect 108 4523 117 4557
rect 117 4523 160 4557
rect 1766 4523 1818 4557
rect 5082 4523 5134 4557
rect 10056 4523 10099 4557
rect 10099 4523 10108 4557
rect 108 4514 160 4523
rect 1766 4514 1818 4523
rect 5082 4514 5134 4523
rect 10056 4514 10108 4523
rect -509 4343 -457 4395
rect 10427 4406 10479 4415
rect 10427 4288 10436 4406
rect 10436 4288 10470 4406
rect 10470 4288 10479 4406
rect 10427 4279 10479 4288
rect -638 4120 -586 4172
rect -380 4132 -328 4184
rect 108 4168 160 4177
rect 1766 4168 1818 4177
rect 5082 4168 5134 4177
rect 8398 4168 8450 4177
rect 10056 4168 10108 4177
rect 108 4134 117 4168
rect 117 4134 160 4168
rect 1766 4134 1818 4168
rect 5082 4134 5134 4168
rect 8398 4134 8450 4168
rect 10056 4134 10099 4168
rect 10099 4134 10108 4168
rect 108 4125 160 4134
rect 1766 4125 1818 4134
rect 5082 4125 5134 4134
rect 8398 4125 8450 4134
rect 10056 4125 10108 4134
rect -509 3987 -457 4039
rect -380 3900 -328 3952
rect -638 3764 -586 3816
rect -509 3631 -457 3683
rect -380 3544 -327 3596
rect -638 3408 -586 3460
rect 108 3894 160 3946
rect 1766 3894 1818 3946
rect 3424 3894 3476 3946
rect 5082 3894 5134 3946
rect 6740 3894 6792 3947
rect 8398 3894 8450 3946
rect 10056 3894 10108 3946
rect 108 3538 160 3590
rect 1766 3538 1818 3590
rect 3424 3538 3476 3590
rect 5082 3538 5134 3590
rect 8398 3538 8450 3590
rect 10056 3538 10108 3590
rect 6740 3414 6792 3466
rect 10649 4867 10701 4919
rect 10780 4688 10832 4740
rect 10649 4511 10701 4563
rect 10780 4332 10832 4384
rect 10951 4406 11003 4415
rect 10951 4288 10960 4406
rect 10960 4288 10994 4406
rect 10994 4288 11003 4406
rect 10951 4279 11003 4288
rect 10649 4155 10701 4207
rect 10780 3976 10832 4028
rect 10649 3799 10701 3851
rect 10545 3676 10597 3728
rect 10780 3620 10832 3672
rect 10551 3556 10603 3608
rect 10651 3442 10703 3494
rect 108 3288 160 3297
rect 1766 3288 1818 3297
rect 5082 3288 5134 3297
rect 8398 3288 8450 3297
rect 10056 3288 10108 3297
rect 108 3254 117 3288
rect 117 3254 160 3288
rect 1766 3254 1818 3288
rect 5082 3254 5134 3288
rect 8398 3254 8450 3288
rect 10056 3254 10099 3288
rect 10099 3254 10108 3288
rect 108 3245 160 3254
rect 1766 3245 1818 3254
rect 5082 3245 5134 3254
rect 8398 3245 8450 3254
rect 10056 3245 10108 3254
rect 10780 3264 10832 3316
rect 1462 2549 1514 2558
rect 5236 2549 5288 2558
rect 8702 2549 8754 2558
rect 1462 2515 1514 2549
rect 5236 2515 5288 2549
rect 8702 2515 8754 2549
rect 1462 2506 1514 2515
rect 5236 2506 5288 2515
rect 8702 2506 8754 2515
rect 3424 2105 3476 2114
rect 3424 2071 3433 2105
rect 3433 2071 3467 2105
rect 3467 2071 3476 2105
rect 3424 2062 3476 2071
rect 6740 2105 6792 2114
rect 6740 2071 6749 2105
rect 6749 2071 6783 2105
rect 6783 2071 6792 2105
rect 6740 2062 6792 2071
rect 3144 1924 3196 1976
rect 4731 1924 4783 1976
rect 6963 1924 7015 1976
rect 108 1827 160 1879
rect 1766 1827 1818 1879
rect 3424 1827 3476 1879
rect 5082 1827 5134 1879
rect 6740 1827 6792 1879
rect 8398 1827 8450 1879
rect 10056 1827 10108 1879
rect 3144 1684 3196 1736
rect 4731 1684 4783 1736
rect 6963 1684 7015 1736
rect 108 1587 160 1639
rect 1766 1587 1818 1639
rect 3424 1587 3476 1639
rect 5082 1587 5134 1639
rect 6740 1587 6792 1639
rect 8398 1587 8450 1639
rect 10056 1587 10108 1639
rect 3144 1444 3196 1496
rect 4731 1444 4783 1496
rect 6963 1444 7015 1496
rect 108 1347 160 1399
rect 1766 1347 1818 1399
rect 3424 1347 3476 1399
rect 5082 1347 5134 1399
rect 6740 1347 6792 1399
rect 8398 1347 8450 1399
rect 10056 1347 10108 1399
rect 3144 1204 3196 1256
rect 4731 1204 4783 1256
rect 6963 1204 7015 1256
rect 108 1107 160 1159
rect 1766 1107 1818 1159
rect 3424 1107 3476 1159
rect 5082 1107 5134 1159
rect 6740 1107 6792 1159
rect 8398 1107 8450 1159
rect 10056 1107 10108 1159
rect 3144 964 3196 1016
rect 4731 964 4783 1016
rect 6963 964 7015 1016
rect 108 867 160 919
rect 1766 867 1818 919
rect 3424 867 3476 919
rect 5082 867 5134 919
rect 6740 867 6792 919
rect 8398 867 8450 919
rect 10056 867 10108 919
rect 3144 724 3196 776
rect 4731 724 4783 776
rect 6963 724 7015 776
rect 108 627 160 679
rect 1766 627 1818 679
rect 3424 627 3476 679
rect 5082 627 5134 679
rect 6740 627 6792 679
rect 8398 627 8450 679
rect 10056 627 10108 679
rect 3144 484 3196 536
rect 4731 484 4783 536
rect 6963 484 7015 536
rect 108 387 160 439
rect 1766 387 1818 439
rect 3424 387 3476 439
rect 5082 387 5134 439
rect 6740 387 6792 439
rect 8398 387 8450 439
rect 10056 387 10108 439
rect 3144 244 3196 296
rect 4731 244 4783 296
rect 6963 244 7015 296
rect 108 147 160 199
rect 1766 147 1818 199
rect 3424 147 3476 199
rect 5082 147 5134 199
rect 6740 147 6792 199
rect 8398 147 8450 199
rect 10056 147 10108 199
rect 3424 17 3476 26
rect 3424 -17 3433 17
rect 3433 -17 3467 17
rect 3467 -17 3476 17
rect 3424 -26 3476 -17
rect 6740 16 6792 25
rect 6740 -18 6749 16
rect 6749 -18 6783 16
rect 6783 -18 6792 16
rect 6740 -27 6792 -18
rect 1462 -427 1514 -418
rect 5236 -427 5288 -418
rect 8702 -427 8754 -418
rect 1462 -461 1514 -427
rect 5236 -461 5288 -427
rect 8702 -461 8754 -427
rect 1462 -470 1514 -461
rect 5236 -470 5288 -461
rect 8702 -470 8754 -461
<< metal2 >>
rect -619 7855 -545 7864
rect -619 7725 -610 7855
rect -554 7725 -545 7855
rect -619 7716 -545 7725
rect 97 7855 171 7864
rect 97 7725 106 7855
rect 162 7725 171 7855
rect 97 7716 171 7725
rect 1755 7855 1829 7864
rect 1755 7725 1764 7855
rect 1820 7725 1829 7855
rect 1755 7716 1829 7725
rect 5071 7855 5145 7864
rect 5071 7725 5080 7855
rect 5136 7725 5145 7855
rect 5071 7716 5145 7725
rect 8387 7855 8461 7864
rect 8387 7725 8396 7855
rect 8452 7725 8461 7855
rect 8387 7716 8461 7725
rect 10045 7855 10119 7864
rect 10045 7725 10054 7855
rect 10110 7725 10119 7855
rect 10045 7716 10119 7725
rect 10734 7855 10808 7864
rect 10734 7725 10743 7855
rect 10799 7725 10808 7855
rect 10734 7716 10808 7725
rect -614 7223 -550 7716
rect 102 7510 166 7716
rect 102 7458 108 7510
rect 160 7458 166 7510
rect 102 7336 166 7458
rect 102 7284 108 7336
rect 160 7284 166 7336
rect -614 7171 -608 7223
rect -556 7171 -550 7223
rect -614 6858 -550 7171
rect -361 7225 -287 7234
rect -361 7169 -352 7225
rect -296 7169 -287 7225
rect -361 7160 -287 7169
rect -614 6806 -608 6858
rect -556 6806 -550 6858
rect -614 6493 -550 6806
rect -614 6441 -608 6493
rect -556 6441 -550 6493
rect -614 6435 -550 6441
rect -485 7115 -421 7121
rect -485 7063 -479 7115
rect -427 7063 -421 7115
rect -485 6750 -421 7063
rect 102 7087 166 7284
rect 102 7035 108 7087
rect 160 7035 166 7087
rect -361 6860 -287 6869
rect -361 6804 -352 6860
rect -296 6804 -287 6860
rect -361 6795 -287 6804
rect 102 6838 166 7035
rect -485 6698 -479 6750
rect -427 6698 -421 6750
rect -485 6385 -421 6698
rect 102 6786 108 6838
rect 160 6786 166 6838
rect 102 6589 166 6786
rect 102 6537 108 6589
rect 160 6537 166 6589
rect -356 6481 -141 6487
rect -356 6429 -350 6481
rect -298 6429 -141 6481
rect -356 6423 -141 6429
rect -485 6369 -479 6385
rect -765 6333 -479 6369
rect -427 6333 -421 6385
rect -765 6305 -421 6333
rect -765 4757 -701 6305
rect -205 6246 -141 6423
rect -485 6182 -141 6246
rect -614 6116 -550 6122
rect -614 6064 -608 6116
rect -556 6064 -550 6116
rect -614 5359 -550 6064
rect -485 6020 -421 6182
rect -485 5968 -479 6020
rect -427 5968 -421 6020
rect -485 5962 -421 5968
rect -356 6116 -292 6122
rect -356 6064 -350 6116
rect -298 6064 -292 6116
rect -624 5350 -550 5359
rect -624 5349 -615 5350
rect -644 5294 -615 5349
rect -559 5294 -550 5350
rect -356 5349 -292 6064
rect -644 5285 -550 5294
rect -386 5285 -292 5349
rect -644 5020 -580 5285
rect -644 4968 -638 5020
rect -586 4968 -580 5020
rect -644 4962 -580 4968
rect -515 5107 -451 5113
rect -515 5055 -509 5107
rect -457 5055 -451 5107
rect -515 4757 -451 5055
rect -386 5031 -322 5285
rect -391 5022 -317 5031
rect -391 4966 -382 5022
rect -326 4966 -317 5022
rect -391 4957 -317 4966
rect -205 4877 -141 6182
rect 102 6340 166 6537
rect 102 6288 108 6340
rect 160 6288 166 6340
rect 102 6091 166 6288
rect 102 6039 108 6091
rect 160 6039 166 6091
rect 102 5842 166 6039
rect 102 5790 108 5842
rect 160 5790 166 5842
rect 102 5593 166 5790
rect 102 5541 108 5593
rect 160 5541 166 5593
rect 102 5344 166 5541
rect 102 5292 108 5344
rect 160 5292 166 5344
rect 102 5100 166 5292
rect 102 5048 108 5100
rect 160 5048 166 5100
rect -107 5015 -33 5024
rect -107 4959 -98 5015
rect -42 4959 -33 5015
rect -107 4950 -33 4959
rect -765 4751 -451 4757
rect -765 4699 -561 4751
rect -509 4699 -451 4751
rect -765 4693 -451 4699
rect -322 4813 -141 4877
rect -322 4670 -258 4813
rect -386 4664 -258 4670
rect -386 4612 -380 4664
rect -328 4612 -258 4664
rect -386 4606 -258 4612
rect -644 4528 -580 4534
rect -644 4476 -638 4528
rect -586 4476 -580 4528
rect -644 4347 -580 4476
rect -386 4445 -322 4606
rect -515 4395 -322 4445
rect -649 4338 -575 4347
rect -649 4282 -640 4338
rect -584 4282 -575 4338
rect -649 4273 -575 4282
rect -515 4343 -509 4395
rect -457 4381 -322 4395
rect -457 4343 -451 4381
rect -644 4172 -580 4273
rect -644 4120 -638 4172
rect -586 4120 -580 4172
rect -644 3816 -580 4120
rect -644 3764 -638 3816
rect -586 3764 -580 3816
rect -644 3460 -580 3764
rect -515 4039 -451 4343
rect -393 4184 -319 4193
rect -100 4187 -40 4950
rect 102 4937 166 5048
rect 102 4885 108 4937
rect 160 4885 166 4937
rect 102 4566 166 4885
rect 102 4514 108 4566
rect 160 4514 166 4566
rect 102 4508 166 4514
rect 1760 7510 1824 7716
rect 1760 7458 1766 7510
rect 1818 7458 1824 7510
rect 1760 7336 1824 7458
rect 5076 7510 5140 7716
rect 5076 7458 5082 7510
rect 5134 7458 5140 7510
rect 1760 7284 1766 7336
rect 1818 7284 1824 7336
rect 1760 7087 1824 7284
rect 3418 7336 3482 7342
rect 3418 7284 3424 7336
rect 3476 7284 3482 7336
rect 3418 7228 3482 7284
rect 5076 7336 5140 7458
rect 8392 7510 8456 7716
rect 8392 7458 8398 7510
rect 8450 7458 8456 7510
rect 5076 7284 5082 7336
rect 5134 7284 5140 7336
rect 3409 7219 3483 7228
rect 3409 7163 3418 7219
rect 3474 7163 3483 7219
rect 3409 7154 3483 7163
rect 1760 7035 1766 7087
rect 1818 7035 1824 7087
rect 1760 6838 1824 7035
rect 1760 6786 1766 6838
rect 1818 6786 1824 6838
rect 1760 6589 1824 6786
rect 1760 6537 1766 6589
rect 1818 6537 1824 6589
rect 1760 6340 1824 6537
rect 1760 6288 1766 6340
rect 1818 6288 1824 6340
rect 1760 6091 1824 6288
rect 1760 6039 1766 6091
rect 1818 6039 1824 6091
rect 1760 5842 1824 6039
rect 1760 5790 1766 5842
rect 1818 5790 1824 5842
rect 1760 5593 1824 5790
rect 1760 5541 1766 5593
rect 1818 5541 1824 5593
rect 1760 5344 1824 5541
rect 1760 5292 1766 5344
rect 1818 5292 1824 5344
rect 1760 5100 1824 5292
rect 1760 5048 1766 5100
rect 1818 5048 1824 5100
rect 1760 4937 1824 5048
rect 3418 7087 3482 7154
rect 3418 7035 3424 7087
rect 3476 7035 3482 7087
rect 3418 6838 3482 7035
rect 3418 6786 3424 6838
rect 3476 6786 3482 6838
rect 3418 6589 3482 6786
rect 3418 6537 3424 6589
rect 3476 6537 3482 6589
rect 3418 6340 3482 6537
rect 3418 6288 3424 6340
rect 3476 6288 3482 6340
rect 3418 6091 3482 6288
rect 5076 7087 5140 7284
rect 5076 7035 5082 7087
rect 5134 7035 5140 7087
rect 5076 6838 5140 7035
rect 6734 7336 6798 7342
rect 6734 7284 6740 7336
rect 6792 7284 6798 7336
rect 6734 7087 6798 7284
rect 6734 7035 6740 7087
rect 6792 7035 6798 7087
rect 6734 6865 6798 7035
rect 8392 7336 8456 7458
rect 8392 7284 8398 7336
rect 8450 7284 8456 7336
rect 8392 7087 8456 7284
rect 8392 7035 8398 7087
rect 8450 7035 8456 7087
rect 5076 6786 5082 6838
rect 5134 6786 5140 6838
rect 6725 6856 6799 6865
rect 6725 6800 6734 6856
rect 6790 6838 6799 6856
rect 6725 6791 6740 6800
rect 5076 6589 5140 6786
rect 5076 6537 5082 6589
rect 5134 6537 5140 6589
rect 5076 6340 5140 6537
rect 5076 6288 5082 6340
rect 5134 6288 5140 6340
rect 3418 6039 3424 6091
rect 3476 6039 3482 6091
rect 3418 5842 3482 6039
rect 3418 5790 3424 5842
rect 3476 5790 3482 5842
rect 3418 5593 3482 5790
rect 3418 5541 3424 5593
rect 3476 5541 3482 5593
rect 3418 5344 3482 5541
rect 3418 5292 3424 5344
rect 3476 5292 3482 5344
rect 3418 5075 3482 5292
rect 4300 6234 4364 6240
rect 4300 6182 4306 6234
rect 4358 6182 4364 6234
rect 4300 5985 4364 6182
rect 4300 5933 4306 5985
rect 4358 5933 4364 5985
rect 4300 5736 4364 5933
rect 4300 5684 4306 5736
rect 4358 5684 4364 5736
rect 4300 5487 4364 5684
rect 4300 5435 4306 5487
rect 4358 5435 4364 5487
rect 4300 5238 4364 5435
rect 4300 5186 4306 5238
rect 4358 5186 4364 5238
rect 3418 5011 3678 5075
rect 1760 4885 1766 4937
rect 1818 4885 1824 4937
rect 1760 4566 1824 4885
rect 3418 4807 3482 4813
rect 3418 4755 3424 4807
rect 3476 4755 3482 4807
rect 3418 4749 3482 4755
rect 1760 4514 1766 4566
rect 1818 4514 1824 4566
rect 97 4409 171 4420
rect 1760 4415 1824 4514
rect 97 4281 106 4409
rect 162 4281 171 4409
rect 97 4272 171 4281
rect 1456 4351 1824 4415
rect -393 4128 -384 4184
rect -328 4128 -319 4184
rect -393 4119 -319 4128
rect -109 4178 -35 4187
rect -109 4122 -100 4178
rect -44 4122 -35 4178
rect -109 4113 -35 4122
rect 102 4177 166 4272
rect 102 4125 108 4177
rect 160 4125 166 4177
rect -515 3987 -509 4039
rect -457 3987 -451 4039
rect -515 3683 -451 3987
rect -395 3952 -321 3960
rect -395 3951 -380 3952
rect -395 3895 -386 3951
rect -328 3900 -321 3952
rect -330 3895 -321 3900
rect -395 3886 -321 3895
rect -515 3631 -509 3683
rect -457 3631 -451 3683
rect -515 3625 -451 3631
rect -100 3603 -40 4113
rect 102 3946 166 4125
rect 102 3894 108 3946
rect 160 3894 166 3946
rect -395 3596 -321 3603
rect -395 3594 -380 3596
rect -395 3538 -386 3594
rect -327 3544 -321 3596
rect -330 3538 -321 3544
rect -395 3529 -321 3538
rect -109 3594 -35 3603
rect -109 3538 -100 3594
rect -44 3538 -35 3594
rect -109 3529 -35 3538
rect 102 3590 166 3894
rect 102 3538 108 3590
rect 160 3538 166 3590
rect -644 3408 -638 3460
rect -586 3408 -580 3460
rect -644 3402 -580 3408
rect 102 3297 166 3538
rect 102 3245 108 3297
rect 160 3245 166 3297
rect 102 1879 166 3245
rect 102 1827 108 1879
rect 160 1827 166 1879
rect 102 1639 166 1827
rect 102 1587 108 1639
rect 160 1587 166 1639
rect 102 1399 166 1587
rect 102 1347 108 1399
rect 160 1347 166 1399
rect 102 1159 166 1347
rect 102 1107 108 1159
rect 160 1107 166 1159
rect 102 919 166 1107
rect 102 867 108 919
rect 160 867 166 919
rect 102 679 166 867
rect 102 627 108 679
rect 160 627 166 679
rect 102 439 166 627
rect 102 387 108 439
rect 160 387 166 439
rect 102 199 166 387
rect 102 147 108 199
rect 160 147 166 199
rect 102 -77 166 147
rect 1456 2558 1520 4351
rect 1760 4177 1824 4183
rect 1760 4125 1766 4177
rect 1818 4125 1824 4177
rect 1760 3946 1824 4125
rect 3424 3953 3476 4749
rect 1760 3894 1766 3946
rect 1818 3894 1824 3946
rect 1760 3590 1824 3894
rect 3409 3946 3483 3953
rect 3409 3944 3424 3946
rect 3409 3888 3418 3944
rect 3476 3894 3483 3946
rect 3474 3888 3483 3894
rect 3409 3879 3483 3888
rect 1760 3538 1766 3590
rect 1818 3538 1824 3590
rect 1760 3297 1824 3538
rect 3409 3590 3483 3597
rect 3409 3588 3424 3590
rect 3409 3532 3418 3588
rect 3476 3538 3483 3590
rect 3474 3532 3483 3538
rect 3409 3523 3483 3532
rect 1760 3245 1766 3297
rect 1818 3245 1824 3297
rect 1760 3239 1824 3245
rect 3133 2915 3207 2924
rect 3133 2859 3142 2915
rect 3198 2859 3207 2915
rect 3133 2850 3207 2859
rect 1456 2506 1462 2558
rect 1514 2506 1520 2558
rect 97 -86 171 -77
rect 97 -216 106 -86
rect 162 -216 171 -86
rect 97 -225 171 -216
rect 1456 -418 1520 2506
rect 1755 2315 1829 2324
rect 1755 2259 1764 2315
rect 1820 2259 1829 2315
rect 1755 2250 1829 2259
rect 1766 1879 1818 2250
rect 3144 1982 3196 2850
rect 3614 2724 3678 5011
rect 4300 4705 4364 5186
rect 4300 4653 4306 4705
rect 4358 4653 4364 4705
rect 3609 2715 3683 2724
rect 3609 2659 3618 2715
rect 3674 2659 3683 2715
rect 3609 2650 3683 2659
rect 3413 2515 3487 2524
rect 3413 2459 3422 2515
rect 3478 2459 3487 2515
rect 3413 2450 3487 2459
rect 3424 2120 3476 2450
rect 4300 2324 4364 4653
rect 5076 6091 5140 6288
rect 6734 6786 6740 6791
rect 6792 6791 6799 6838
rect 8392 6838 8456 7035
rect 6792 6786 6798 6791
rect 6734 6589 6798 6786
rect 6734 6537 6740 6589
rect 6792 6537 6798 6589
rect 6734 6340 6798 6537
rect 6734 6288 6740 6340
rect 6792 6288 6798 6340
rect 5076 6039 5082 6091
rect 5134 6039 5140 6091
rect 5076 5842 5140 6039
rect 5076 5790 5082 5842
rect 5134 5790 5140 5842
rect 5076 5593 5140 5790
rect 5076 5541 5082 5593
rect 5134 5541 5140 5593
rect 5076 5344 5140 5541
rect 5076 5292 5082 5344
rect 5134 5292 5140 5344
rect 5076 5100 5140 5292
rect 5076 5048 5082 5100
rect 5134 5048 5140 5100
rect 5076 4937 5140 5048
rect 5076 4885 5082 4937
rect 5134 4885 5140 4937
rect 5076 4572 5140 4885
rect 5956 6234 6020 6240
rect 5956 6182 5962 6234
rect 6014 6182 6020 6234
rect 5956 5985 6020 6182
rect 5956 5933 5962 5985
rect 6014 5933 6020 5985
rect 5956 5736 6020 5933
rect 5956 5684 5962 5736
rect 6014 5684 6020 5736
rect 5956 5487 6020 5684
rect 5956 5435 5962 5487
rect 6014 5435 6020 5487
rect 5956 5238 6020 5435
rect 5956 5186 5962 5238
rect 6014 5186 6020 5238
rect 5956 4705 6020 5186
rect 6734 6091 6798 6288
rect 6734 6039 6740 6091
rect 6792 6039 6798 6091
rect 6734 5842 6798 6039
rect 6734 5790 6740 5842
rect 6792 5790 6798 5842
rect 6734 5593 6798 5790
rect 6734 5541 6740 5593
rect 6792 5541 6798 5593
rect 6734 5344 6798 5541
rect 6734 5292 6740 5344
rect 6792 5292 6798 5344
rect 6734 5075 6798 5292
rect 5956 4653 5962 4705
rect 6014 4653 6020 4705
rect 5076 4566 5294 4572
rect 5076 4514 5082 4566
rect 5134 4514 5294 4566
rect 5076 4508 5294 4514
rect 5071 4410 5145 4421
rect 5071 4282 5080 4410
rect 5136 4282 5145 4410
rect 5071 4273 5145 4282
rect 5076 4177 5140 4273
rect 5076 4125 5082 4177
rect 5134 4125 5140 4177
rect 5076 3946 5140 4125
rect 5076 3894 5082 3946
rect 5134 3894 5140 3946
rect 5076 3590 5140 3894
rect 5076 3538 5082 3590
rect 5134 3538 5140 3590
rect 5076 3297 5140 3538
rect 5076 3245 5082 3297
rect 5134 3245 5140 3297
rect 5076 3239 5140 3245
rect 4720 3115 4794 3124
rect 4720 3059 4729 3115
rect 4785 3059 4794 3115
rect 4720 3050 4794 3059
rect 4295 2315 4369 2324
rect 4295 2259 4304 2315
rect 4360 2259 4369 2315
rect 4295 2250 4369 2259
rect 3418 2114 3482 2120
rect 3418 2062 3424 2114
rect 3476 2062 3482 2114
rect 3418 2056 3482 2062
rect 3138 1976 3202 1982
rect 3138 1924 3144 1976
rect 3196 1924 3202 1976
rect 3138 1918 3202 1924
rect 1766 1821 1818 1827
rect 3144 1742 3196 1918
rect 3424 1879 3476 2056
rect 4731 1982 4783 3050
rect 5071 2715 5145 2724
rect 5071 2659 5080 2715
rect 5136 2659 5145 2715
rect 5071 2650 5145 2659
rect 4725 1976 4789 1982
rect 4725 1924 4731 1976
rect 4783 1924 4789 1976
rect 4725 1918 4789 1924
rect 3424 1821 3476 1827
rect 4731 1742 4783 1918
rect 5082 1879 5134 2650
rect 5082 1821 5134 1827
rect 5230 2558 5294 4508
rect 5956 2721 6020 4653
rect 6538 5011 6798 5075
rect 8392 6786 8398 6838
rect 8450 6786 8456 6838
rect 8392 6589 8456 6786
rect 8392 6537 8398 6589
rect 8450 6537 8456 6589
rect 8392 6340 8456 6537
rect 8392 6288 8398 6340
rect 8450 6288 8456 6340
rect 8392 6091 8456 6288
rect 8392 6039 8398 6091
rect 8450 6039 8456 6091
rect 8392 5842 8456 6039
rect 8392 5790 8398 5842
rect 8450 5790 8456 5842
rect 8392 5593 8456 5790
rect 8392 5541 8398 5593
rect 8450 5541 8456 5593
rect 8392 5344 8456 5541
rect 8392 5292 8398 5344
rect 8450 5292 8456 5344
rect 8392 5100 8456 5292
rect 8392 5048 8398 5100
rect 8450 5048 8456 5100
rect 5950 2712 6024 2721
rect 5950 2656 5959 2712
rect 6015 2656 6024 2712
rect 5950 2647 6024 2656
rect 5230 2506 5236 2558
rect 5288 2506 5294 2558
rect 3138 1736 3202 1742
rect 3138 1684 3144 1736
rect 3196 1684 3202 1736
rect 3138 1678 3202 1684
rect 4725 1736 4789 1742
rect 4725 1684 4731 1736
rect 4783 1684 4789 1736
rect 4725 1678 4789 1684
rect 1766 1639 1818 1645
rect 1766 1581 1818 1587
rect 3144 1502 3196 1678
rect 3424 1639 3476 1645
rect 3424 1581 3476 1587
rect 4731 1502 4783 1678
rect 5082 1639 5134 1645
rect 5082 1581 5134 1587
rect 3138 1496 3202 1502
rect 3138 1444 3144 1496
rect 3196 1444 3202 1496
rect 3138 1438 3202 1444
rect 4725 1496 4789 1502
rect 4725 1444 4731 1496
rect 4783 1444 4789 1496
rect 4725 1438 4789 1444
rect 1766 1399 1818 1405
rect 1766 1341 1818 1347
rect 3144 1262 3196 1438
rect 3424 1399 3476 1405
rect 3424 1341 3476 1347
rect 4731 1262 4783 1438
rect 5082 1399 5134 1405
rect 5082 1341 5134 1347
rect 3138 1256 3202 1262
rect 3138 1204 3144 1256
rect 3196 1204 3202 1256
rect 3138 1198 3202 1204
rect 4725 1256 4789 1262
rect 4725 1204 4731 1256
rect 4783 1204 4789 1256
rect 4725 1198 4789 1204
rect 1766 1159 1818 1165
rect 1766 1101 1818 1107
rect 3144 1022 3196 1198
rect 3424 1159 3476 1165
rect 3424 1101 3476 1107
rect 4731 1022 4783 1198
rect 5082 1159 5134 1165
rect 5082 1101 5134 1107
rect 3138 1016 3202 1022
rect 3138 964 3144 1016
rect 3196 964 3202 1016
rect 3138 958 3202 964
rect 4725 1016 4789 1022
rect 4725 964 4731 1016
rect 4783 964 4789 1016
rect 4725 958 4789 964
rect 1766 919 1818 925
rect 1766 861 1818 867
rect 3144 782 3196 958
rect 3424 919 3476 925
rect 3424 861 3476 867
rect 4731 782 4783 958
rect 5082 919 5134 925
rect 5082 861 5134 867
rect 3138 776 3202 782
rect 3138 724 3144 776
rect 3196 724 3202 776
rect 3138 718 3202 724
rect 4725 776 4789 782
rect 4725 724 4731 776
rect 4783 724 4789 776
rect 4725 718 4789 724
rect 1766 679 1818 685
rect 1766 621 1818 627
rect 3144 542 3196 718
rect 3424 679 3476 685
rect 3424 621 3476 627
rect 4731 542 4783 718
rect 5082 679 5134 685
rect 5082 621 5134 627
rect 3138 536 3202 542
rect 3138 484 3144 536
rect 3196 484 3202 536
rect 3138 478 3202 484
rect 4725 536 4789 542
rect 4725 484 4731 536
rect 4783 484 4789 536
rect 4725 478 4789 484
rect 1766 439 1818 445
rect 1766 381 1818 387
rect 3144 302 3196 478
rect 3424 439 3476 445
rect 3424 381 3476 387
rect 4731 302 4783 478
rect 5082 439 5134 445
rect 5082 381 5134 387
rect 3138 296 3202 302
rect 3138 244 3144 296
rect 3196 244 3202 296
rect 3138 238 3202 244
rect 4725 296 4789 302
rect 4725 244 4731 296
rect 4783 244 4789 296
rect 4725 238 4789 244
rect 1766 199 1818 205
rect 1766 141 1818 147
rect 3424 199 3476 205
rect 3424 32 3476 147
rect 5082 199 5134 205
rect 5082 141 5134 147
rect 3418 26 3482 32
rect 3418 -26 3424 26
rect 3476 -26 3482 26
rect 3418 -32 3482 -26
rect 1456 -470 1462 -418
rect 1514 -470 1520 -418
rect 1456 -476 1520 -470
rect 5230 -418 5294 2506
rect 6538 2324 6602 5011
rect 8392 4937 8456 5048
rect 8392 4885 8398 4937
rect 8450 4885 8456 4937
rect 6734 4807 6798 4813
rect 6734 4755 6740 4807
rect 6792 4755 6798 4807
rect 6734 4749 6798 4755
rect 6740 3954 6792 4749
rect 8392 4415 8456 4885
rect 10050 7510 10114 7716
rect 10050 7458 10056 7510
rect 10108 7458 10114 7510
rect 10050 7336 10114 7458
rect 10050 7284 10056 7336
rect 10108 7284 10114 7336
rect 10050 7087 10114 7284
rect 10739 7510 10803 7716
rect 10739 7458 10745 7510
rect 10797 7458 10803 7510
rect 10739 7376 10803 7458
rect 10739 7324 10745 7376
rect 10797 7324 10803 7376
rect 10050 7035 10056 7087
rect 10108 7035 10114 7087
rect 10050 6838 10114 7035
rect 10050 6786 10056 6838
rect 10108 6786 10114 6838
rect 10050 6589 10114 6786
rect 10050 6537 10056 6589
rect 10108 6537 10114 6589
rect 10050 6340 10114 6537
rect 10050 6288 10056 6340
rect 10108 6288 10114 6340
rect 10050 6091 10114 6288
rect 10609 7198 10673 7204
rect 10609 7146 10615 7198
rect 10667 7146 10673 7198
rect 10609 6842 10673 7146
rect 10609 6790 10615 6842
rect 10667 6790 10673 6842
rect 10609 6486 10673 6790
rect 10609 6434 10615 6486
rect 10667 6434 10673 6486
rect 10609 6142 10673 6434
rect 10739 7020 10803 7324
rect 10739 6968 10745 7020
rect 10797 6968 10803 7020
rect 10739 6664 10803 6968
rect 10739 6612 10745 6664
rect 10797 6612 10803 6664
rect 10739 6308 10803 6612
rect 10739 6256 10745 6308
rect 10797 6256 10803 6308
rect 10050 6039 10056 6091
rect 10108 6039 10114 6091
rect 10050 5842 10114 6039
rect 10050 5790 10056 5842
rect 10108 5790 10114 5842
rect 10050 5593 10114 5790
rect 10050 5541 10056 5593
rect 10108 5541 10114 5593
rect 10050 5344 10114 5541
rect 10050 5292 10056 5344
rect 10108 5292 10114 5344
rect 10050 5100 10114 5292
rect 10050 5048 10056 5100
rect 10108 5048 10114 5100
rect 10050 4937 10114 5048
rect 10050 4885 10056 4937
rect 10108 4885 10114 4937
rect 10186 6130 10260 6139
rect 10186 6074 10195 6130
rect 10251 6074 10260 6130
rect 10186 6065 10260 6074
rect 10602 6133 10676 6142
rect 10602 6077 10611 6133
rect 10667 6077 10676 6133
rect 10602 6068 10676 6077
rect 10186 4922 10242 6065
rect 10506 6007 10570 6013
rect 10506 5955 10512 6007
rect 10564 5995 10570 6007
rect 10564 5955 10665 5995
rect 10506 5949 10665 5955
rect 10609 5780 10665 5949
rect 10739 5952 10803 6256
rect 10739 5900 10745 5952
rect 10797 5900 10803 5952
rect 10609 5774 10673 5780
rect 10609 5722 10615 5774
rect 10667 5722 10673 5774
rect 10609 5716 10673 5722
rect 10508 5661 10572 5667
rect 10508 5656 10514 5661
rect 10312 5609 10514 5656
rect 10566 5609 10572 5661
rect 10312 5603 10572 5609
rect 10050 4566 10114 4885
rect 10174 4913 10248 4922
rect 10174 4857 10183 4913
rect 10239 4857 10248 4913
rect 10174 4848 10248 4857
rect 10050 4514 10056 4566
rect 10108 4514 10114 4566
rect 10050 4508 10114 4514
rect 8392 4351 8760 4415
rect 8392 4177 8456 4183
rect 8392 4125 8398 4177
rect 8450 4125 8456 4177
rect 6724 3947 6798 3954
rect 6724 3945 6740 3947
rect 6724 3889 6733 3945
rect 6792 3894 6798 3947
rect 6789 3889 6798 3894
rect 6724 3880 6798 3889
rect 8392 3946 8456 4125
rect 8392 3894 8398 3946
rect 8450 3894 8456 3946
rect 8392 3590 8456 3894
rect 8392 3538 8398 3590
rect 8450 3538 8456 3590
rect 6734 3466 6798 3472
rect 6734 3414 6740 3466
rect 6792 3414 6798 3466
rect 6734 3408 6798 3414
rect 6740 2524 6792 3408
rect 8392 3297 8456 3538
rect 8392 3245 8398 3297
rect 8450 3245 8456 3297
rect 8392 3239 8456 3245
rect 6952 2915 7026 2924
rect 6952 2859 6961 2915
rect 7017 2859 7026 2915
rect 6952 2850 7026 2859
rect 6729 2515 6803 2524
rect 6729 2459 6738 2515
rect 6794 2459 6803 2515
rect 6729 2450 6803 2459
rect 6533 2315 6607 2324
rect 6533 2259 6542 2315
rect 6598 2259 6607 2315
rect 6533 2250 6607 2259
rect 6740 2120 6792 2450
rect 6734 2114 6798 2120
rect 6734 2062 6740 2114
rect 6792 2062 6798 2114
rect 6734 2056 6798 2062
rect 6740 1879 6792 2056
rect 6963 1982 7015 2850
rect 8696 2558 8760 4351
rect 10045 4410 10119 4421
rect 10045 4284 10054 4410
rect 10110 4284 10119 4410
rect 10045 4273 10119 4284
rect 8696 2506 8702 2558
rect 8754 2506 8760 2558
rect 8387 2315 8461 2324
rect 8387 2259 8396 2315
rect 8452 2259 8461 2315
rect 8387 2250 8461 2259
rect 6957 1976 7021 1982
rect 6957 1924 6963 1976
rect 7015 1924 7021 1976
rect 6957 1918 7021 1924
rect 6740 1821 6792 1827
rect 6963 1742 7015 1918
rect 8398 1879 8450 2250
rect 8398 1821 8450 1827
rect 6957 1736 7021 1742
rect 6957 1684 6963 1736
rect 7015 1684 7021 1736
rect 6957 1678 7021 1684
rect 6740 1639 6792 1645
rect 6740 1581 6792 1587
rect 6963 1502 7015 1678
rect 8398 1639 8450 1645
rect 8398 1581 8450 1587
rect 6957 1496 7021 1502
rect 6957 1444 6963 1496
rect 7015 1444 7021 1496
rect 6957 1438 7021 1444
rect 6740 1399 6792 1405
rect 6740 1341 6792 1347
rect 6963 1262 7015 1438
rect 8398 1399 8450 1405
rect 8398 1341 8450 1347
rect 6957 1256 7021 1262
rect 6957 1204 6963 1256
rect 7015 1204 7021 1256
rect 6957 1198 7021 1204
rect 6740 1159 6792 1165
rect 6740 1101 6792 1107
rect 6963 1022 7015 1198
rect 8398 1159 8450 1165
rect 8398 1101 8450 1107
rect 6957 1016 7021 1022
rect 6957 964 6963 1016
rect 7015 964 7021 1016
rect 6957 958 7021 964
rect 6740 919 6792 925
rect 6740 861 6792 867
rect 6963 782 7015 958
rect 8398 919 8450 925
rect 8398 861 8450 867
rect 6957 776 7021 782
rect 6957 724 6963 776
rect 7015 724 7021 776
rect 6957 718 7021 724
rect 6740 679 6792 685
rect 6740 621 6792 627
rect 6963 542 7015 718
rect 8398 679 8450 685
rect 8398 621 8450 627
rect 6957 536 7021 542
rect 6957 484 6963 536
rect 7015 484 7021 536
rect 6957 478 7021 484
rect 6740 439 6792 445
rect 6740 381 6792 387
rect 6963 302 7015 478
rect 8398 439 8450 445
rect 8398 381 8450 387
rect 6957 296 7021 302
rect 6957 244 6963 296
rect 7015 244 7021 296
rect 6957 238 7021 244
rect 6740 199 6792 205
rect 6740 31 6792 147
rect 8398 199 8450 205
rect 8398 141 8450 147
rect 6734 25 6798 31
rect 6734 -27 6740 25
rect 6792 -27 6798 25
rect 6734 -33 6798 -27
rect 5230 -470 5236 -418
rect 5288 -470 5294 -418
rect 5230 -480 5294 -470
rect 8696 -418 8760 2506
rect 10050 4177 10114 4273
rect 10050 4125 10056 4177
rect 10108 4125 10114 4177
rect 10050 3946 10114 4125
rect 10050 3894 10056 3946
rect 10108 3894 10114 3946
rect 10050 3590 10114 3894
rect 10312 3796 10368 5603
rect 10609 5569 10665 5716
rect 10539 5513 10665 5569
rect 10739 5596 10803 5900
rect 10739 5544 10745 5596
rect 10797 5544 10803 5596
rect 10416 4415 10490 4421
rect 10416 4410 10427 4415
rect 10479 4410 10490 4415
rect 10416 4284 10425 4410
rect 10481 4284 10490 4410
rect 10416 4279 10427 4284
rect 10479 4279 10490 4284
rect 10416 4273 10490 4279
rect 10303 3787 10377 3796
rect 10303 3731 10312 3787
rect 10368 3731 10377 3787
rect 10303 3722 10377 3731
rect 10539 3734 10595 5513
rect 10739 5462 10803 5544
rect 10739 5410 10745 5462
rect 10797 5410 10803 5462
rect 10739 5404 10803 5410
rect 10774 5096 10838 5102
rect 10774 5044 10780 5096
rect 10832 5044 10838 5096
rect 10635 4920 10709 4929
rect 10635 4864 10644 4920
rect 10700 4919 10709 4920
rect 10701 4867 10709 4919
rect 10700 4864 10709 4867
rect 10635 4855 10709 4864
rect 10643 4563 10707 4855
rect 10643 4511 10649 4563
rect 10701 4511 10707 4563
rect 10643 4207 10707 4511
rect 10643 4155 10649 4207
rect 10701 4155 10707 4207
rect 10643 3851 10707 4155
rect 10643 3799 10649 3851
rect 10701 3799 10707 3851
rect 10643 3793 10707 3799
rect 10774 4740 10838 5044
rect 10774 4688 10780 4740
rect 10832 4688 10838 4740
rect 10774 4421 10838 4688
rect 10774 4410 10848 4421
rect 10774 4384 10783 4410
rect 10774 4332 10780 4384
rect 10774 4284 10783 4332
rect 10839 4284 10848 4410
rect 10774 4273 10848 4284
rect 10940 4415 11014 4421
rect 10940 4410 10951 4415
rect 11003 4410 11014 4415
rect 10940 4284 10949 4410
rect 11005 4284 11014 4410
rect 10940 4279 10951 4284
rect 11003 4279 11014 4284
rect 10940 4273 11014 4279
rect 10774 4028 10838 4273
rect 10774 3976 10780 4028
rect 10832 3976 10838 4028
rect 10539 3729 10603 3734
rect 10539 3728 10704 3729
rect 10050 3538 10056 3590
rect 10108 3538 10114 3590
rect 10312 3613 10368 3722
rect 10539 3676 10545 3728
rect 10597 3676 10704 3728
rect 10539 3673 10704 3676
rect 10539 3670 10603 3673
rect 10545 3613 10609 3614
rect 10312 3608 10609 3613
rect 10312 3557 10551 3608
rect 10545 3556 10551 3557
rect 10603 3556 10609 3608
rect 10545 3550 10609 3556
rect 10050 3297 10114 3538
rect 10648 3500 10704 3673
rect 10774 3672 10838 3976
rect 10774 3620 10780 3672
rect 10832 3620 10838 3672
rect 10645 3494 10709 3500
rect 10645 3442 10651 3494
rect 10703 3442 10709 3494
rect 10645 3436 10709 3442
rect 10050 3245 10056 3297
rect 10108 3245 10114 3297
rect 10774 3316 10838 3620
rect 10774 3264 10780 3316
rect 10832 3264 10838 3316
rect 10774 3258 10838 3264
rect 10050 1879 10114 3245
rect 10050 1827 10056 1879
rect 10108 1827 10114 1879
rect 10050 1639 10114 1827
rect 10050 1587 10056 1639
rect 10108 1587 10114 1639
rect 10050 1399 10114 1587
rect 10050 1347 10056 1399
rect 10108 1347 10114 1399
rect 10050 1159 10114 1347
rect 10050 1107 10056 1159
rect 10108 1107 10114 1159
rect 10050 919 10114 1107
rect 10050 867 10056 919
rect 10108 867 10114 919
rect 10050 679 10114 867
rect 10050 627 10056 679
rect 10108 627 10114 679
rect 10050 439 10114 627
rect 10050 387 10056 439
rect 10108 387 10114 439
rect 10050 199 10114 387
rect 10050 147 10056 199
rect 10108 147 10114 199
rect 10050 -77 10114 147
rect 10045 -86 10119 -77
rect 10045 -216 10054 -86
rect 10110 -216 10119 -86
rect 10045 -225 10119 -216
rect 8696 -470 8702 -418
rect 8754 -470 8760 -418
rect 8696 -476 8760 -470
<< via2 >>
rect -610 7725 -554 7855
rect 106 7725 162 7855
rect 1764 7725 1820 7855
rect 5080 7725 5136 7855
rect 8396 7725 8452 7855
rect 10054 7725 10110 7855
rect 10743 7725 10799 7855
rect -352 7223 -296 7225
rect -352 7171 -350 7223
rect -350 7171 -298 7223
rect -298 7171 -296 7223
rect -352 7169 -296 7171
rect -352 6858 -296 6860
rect -352 6806 -350 6858
rect -350 6806 -298 6858
rect -298 6806 -296 6858
rect -352 6804 -296 6806
rect -615 5294 -559 5350
rect -382 5020 -326 5022
rect -382 4968 -380 5020
rect -380 4968 -328 5020
rect -328 4968 -326 5020
rect -382 4966 -326 4968
rect -98 4959 -42 5015
rect -640 4282 -584 4338
rect 3418 7163 3474 7219
rect 6734 6838 6790 6856
rect 6734 6800 6740 6838
rect 6740 6800 6790 6838
rect 106 4281 162 4409
rect -384 4132 -380 4184
rect -380 4132 -328 4184
rect -384 4128 -328 4132
rect -100 4122 -44 4178
rect -386 3900 -380 3951
rect -380 3900 -330 3951
rect -386 3895 -330 3900
rect -386 3544 -380 3594
rect -380 3544 -330 3594
rect -386 3538 -330 3544
rect -100 3538 -44 3594
rect 3418 3894 3424 3944
rect 3424 3894 3474 3944
rect 3418 3888 3474 3894
rect 3418 3538 3424 3588
rect 3424 3538 3474 3588
rect 3418 3532 3474 3538
rect 3142 2859 3198 2915
rect 106 -216 162 -86
rect 1764 2259 1820 2315
rect 3618 2659 3674 2715
rect 3422 2459 3478 2515
rect 5080 4282 5136 4410
rect 4729 3059 4785 3115
rect 4304 2259 4360 2315
rect 5080 2659 5136 2715
rect 5959 2656 6015 2712
rect 10195 6074 10251 6130
rect 10611 6130 10667 6133
rect 10611 6078 10615 6130
rect 10615 6078 10667 6130
rect 10611 6077 10667 6078
rect 10183 4857 10239 4913
rect 6733 3894 6740 3945
rect 6740 3894 6789 3945
rect 6733 3889 6789 3894
rect 6961 2859 7017 2915
rect 6738 2459 6794 2515
rect 6542 2259 6598 2315
rect 10054 4284 10110 4410
rect 8396 2259 8452 2315
rect 10425 4284 10427 4410
rect 10427 4284 10479 4410
rect 10479 4284 10481 4410
rect 10312 3731 10368 3787
rect 10644 4919 10700 4920
rect 10644 4867 10649 4919
rect 10649 4867 10700 4919
rect 10644 4864 10700 4867
rect 10783 4384 10839 4410
rect 10783 4332 10832 4384
rect 10832 4332 10839 4384
rect 10783 4284 10839 4332
rect 10949 4284 10951 4410
rect 10951 4284 11003 4410
rect 11003 4284 11005 4410
rect 10054 -216 10110 -86
<< metal3 >>
rect -619 7855 10808 7864
rect -619 7725 -610 7855
rect -554 7725 106 7855
rect 162 7725 1764 7855
rect 1820 7725 5080 7855
rect 5136 7725 8396 7855
rect 8452 7725 10054 7855
rect 10110 7725 10743 7855
rect 10799 7725 10808 7855
rect -619 7716 10808 7725
rect -361 7225 -287 7234
rect 3409 7225 3483 7228
rect -361 7169 -352 7225
rect -296 7219 3483 7225
rect -296 7169 3418 7219
rect -361 7165 3418 7169
rect -361 7160 -287 7165
rect 3409 7163 3418 7165
rect 3474 7163 3483 7219
rect 3409 7154 3483 7163
rect -361 6861 -287 6869
rect 6725 6861 6799 6865
rect -361 6860 6799 6861
rect -361 6804 -352 6860
rect -296 6856 6799 6860
rect -296 6804 6734 6856
rect -361 6801 6734 6804
rect -361 6795 -287 6801
rect 6725 6800 6734 6801
rect 6790 6800 6799 6856
rect 6725 6791 6799 6800
rect 10186 6132 10260 6139
rect 10602 6133 10676 6142
rect 10602 6132 10611 6133
rect 10186 6130 10611 6132
rect 10186 6074 10195 6130
rect 10251 6077 10611 6130
rect 10667 6077 10676 6133
rect 10251 6074 10676 6077
rect 10186 6072 10676 6074
rect 10186 6065 10260 6072
rect 10602 6068 10676 6072
rect -701 5350 -550 5359
rect -701 5294 -615 5350
rect -559 5294 -550 5350
rect -701 5285 -550 5294
rect -391 5022 -317 5031
rect -391 4966 -382 5022
rect -326 5017 -317 5022
rect -107 5017 -33 5024
rect -326 5015 -33 5017
rect -326 4966 -98 5015
rect -391 4959 -98 4966
rect -42 4959 -33 5015
rect -391 4957 -33 4959
rect -107 4950 -33 4957
rect 10174 4920 10248 4922
rect 10635 4920 10709 4929
rect 10174 4913 10644 4920
rect 10174 4857 10183 4913
rect 10239 4864 10644 4913
rect 10700 4864 10709 4920
rect 10239 4860 10709 4864
rect 10239 4857 10248 4860
rect 10174 4848 10248 4857
rect 10635 4855 10709 4860
rect -649 4420 97 4421
rect 171 4420 11014 4421
rect -649 4410 11014 4420
rect -649 4409 5080 4410
rect -649 4338 106 4409
rect -649 4282 -640 4338
rect -584 4282 106 4338
rect -649 4281 106 4282
rect 162 4282 5080 4409
rect 5136 4284 10054 4410
rect 10110 4284 10425 4410
rect 10481 4284 10783 4410
rect 10839 4284 10949 4410
rect 11005 4284 11014 4410
rect 5136 4282 11014 4284
rect 162 4281 11014 4282
rect -649 4273 11014 4281
rect 97 4272 171 4273
rect -393 4184 -319 4193
rect -393 4128 -384 4184
rect -328 4182 -319 4184
rect -109 4182 -35 4187
rect -328 4178 -35 4182
rect -328 4128 -100 4178
rect -393 4122 -100 4128
rect -44 4122 -35 4178
rect -393 4119 -319 4122
rect -109 4113 -35 4122
rect -395 3951 -321 3960
rect 3409 3951 3483 3953
rect -395 3895 -386 3951
rect -330 3944 3483 3951
rect -330 3895 3418 3944
rect -395 3891 3418 3895
rect -395 3886 -321 3891
rect 3409 3888 3418 3891
rect 3474 3888 3483 3944
rect 3409 3879 3483 3888
rect 6724 3945 6798 3954
rect 6724 3889 6733 3945
rect 6789 3889 6798 3945
rect 6724 3880 6798 3889
rect 6724 3791 6784 3880
rect 10303 3791 10377 3796
rect -356 3787 10377 3791
rect -356 3731 10312 3787
rect 10368 3731 10377 3787
rect -356 3625 -296 3731
rect 10303 3722 10377 3731
rect -395 3594 -296 3625
rect -395 3538 -386 3594
rect -330 3565 -296 3594
rect -109 3594 -35 3603
rect 3409 3594 3483 3597
rect -330 3538 -321 3565
rect -395 3529 -321 3538
rect -109 3538 -100 3594
rect -44 3588 3483 3594
rect -44 3538 3418 3588
rect -109 3534 3418 3538
rect -109 3529 -35 3534
rect 3409 3532 3418 3534
rect 3474 3532 3483 3588
rect 3409 3523 3483 3532
rect 4720 3117 4794 3124
rect 1766 3115 8450 3117
rect 1766 3059 4729 3115
rect 4785 3059 8450 3115
rect 1766 3057 8450 3059
rect 4720 3050 4794 3057
rect 3133 2917 3207 2924
rect 6952 2917 7026 2924
rect 1766 2915 8450 2917
rect 1766 2859 3142 2915
rect 3198 2859 6961 2915
rect 7017 2859 8450 2915
rect 1766 2857 8450 2859
rect 3133 2850 3207 2857
rect 6952 2850 7026 2857
rect 3609 2717 3683 2724
rect 5071 2717 5145 2724
rect 5950 2717 6024 2721
rect 1766 2715 8450 2717
rect 1766 2659 3618 2715
rect 3674 2659 5080 2715
rect 5136 2712 8450 2715
rect 5136 2659 5959 2712
rect 1766 2657 5959 2659
rect 3609 2650 3683 2657
rect 5071 2650 5145 2657
rect 5950 2656 5959 2657
rect 6015 2657 8450 2712
rect 6015 2656 6024 2657
rect 5950 2647 6024 2656
rect 3413 2517 3487 2524
rect 6729 2517 6803 2524
rect 1766 2515 8450 2517
rect 1766 2459 3422 2515
rect 3478 2459 6738 2515
rect 6794 2459 8450 2515
rect 1766 2457 8450 2459
rect 3413 2450 3487 2457
rect 6729 2450 6803 2457
rect 1755 2317 1829 2324
rect 4295 2317 4369 2324
rect 6533 2317 6607 2324
rect 8387 2317 8461 2324
rect 1755 2315 8461 2317
rect 1755 2259 1764 2315
rect 1820 2259 4304 2315
rect 4360 2259 6542 2315
rect 6598 2259 8396 2315
rect 8452 2259 8461 2315
rect 1755 2257 8461 2259
rect 1755 2250 1829 2257
rect 4295 2250 4369 2257
rect 6533 2250 6607 2257
rect 8387 2250 8461 2257
rect 97 -86 10119 -77
rect 97 -216 106 -86
rect 162 -216 10054 -86
rect 10110 -216 10119 -86
rect 97 -225 10119 -216
use sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z  sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z_0
timestamp 1712352531
transform 1 0 -483 0 1 4245
box -328 -1039 328 1039
use sky130_fd_pr__nfet_g5v0d10v5_GLAJGT  sky130_fd_pr__nfet_g5v0d10v5_GLAJGT_1
timestamp 1712352531
transform 1 0 5108 0 1 1044
box -5173 -1109 5173 1109
use sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z  sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z_0
timestamp 1712352531
transform 0 -1 10707 -1 0 4180
box -1089 -327 1089 327
use sky130_fd_pr__nfet_g5v0d10v5_T82T27  sky130_fd_pr__nfet_g5v0d10v5_T82T27_1
timestamp 1712352531
transform 1 0 5108 0 1 3711
box -5173 -505 5173 505
use sky130_fd_pr__pfet_g5v0d10v5_3HV7M9  sky130_fd_pr__pfet_g5v0d10v5_3HV7M9_0
timestamp 1712352531
transform 1 0 5108 0 1 4807
box -5203 -362 5203 362
use sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4  sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4_0
timestamp 1712352531
transform 1 0 -453 0 1 6670
box -358 -909 358 909
use sky130_fd_pr__pfet_g5v0d10v5_8FRRWQ  sky130_fd_pr__pfet_g5v0d10v5_8FRRWQ_0
timestamp 1712352531
transform 1 0 5108 0 1 6279
box -5203 -1300 5203 1300
use sky130_fd_pr__pfet_g5v0d10v5_W8MWAU  sky130_fd_pr__pfet_g5v0d10v5_W8MWAU_0
timestamp 1712352531
transform 0 -1 10673 -1 0 6460
box -1119 -362 1119 362
<< labels >>
rlabel metal2 3424 4230 3424 4230 7 vm
rlabel metal2 3418 3596 3418 3596 7 vn
flabel comment s 995 1104 995 1104 0 FreeSans 1600 0 0 0 dum
flabel comment s 2653 1104 2653 1104 0 FreeSans 1600 0 0 0 Mi0
flabel comment s 4311 1104 4311 1104 0 FreeSans 1600 0 0 0 Mi1
flabel comment s 5969 1104 5969 1104 0 FreeSans 1600 0 0 0 Mi1
flabel comment s 7627 1104 7627 1104 0 FreeSans 1600 0 0 0 Mi0
flabel comment s 9285 1104 9285 1104 0 FreeSans 1600 0 0 0 dum
flabel comment s 9285 3504 9285 3504 0 FreeSans 1600 0 0 0 dum
flabel comment s 7627 3504 7627 3504 0 FreeSans 1600 0 0 0 Mta
flabel comment s 5969 3504 5969 3504 0 FreeSans 1600 0 0 0 Mta
flabel comment s 4311 3504 4311 3504 0 FreeSans 1600 0 0 0 Mb
flabel comment s 2653 3504 2653 3504 0 FreeSans 1600 0 0 0 Mb
flabel comment s 995 3504 995 3504 0 FreeSans 1600 0 0 0 dum
flabel comment s 995 3864 995 3864 0 FreeSans 1600 0 0 0 dum
flabel comment s 2653 3864 2653 3864 0 FreeSans 1600 0 0 0 Mnn0
flabel comment s 4311 3864 4311 3864 0 FreeSans 1600 0 0 0 Mnn0
flabel comment s 5969 3864 5969 3864 0 FreeSans 1600 0 0 0 Mnn1
flabel comment s 7627 3864 7627 3864 0 FreeSans 1600 0 0 0 Mnn1
flabel comment s 9285 3864 9285 3864 0 FreeSans 1600 0 0 0 dum
flabel comment s 9285 4824 9285 4824 0 FreeSans 1600 0 0 0 dum
flabel comment s 7627 4824 7627 4824 0 FreeSans 1600 0 0 0 Mpp1
flabel comment s 5969 4824 5969 4824 0 FreeSans 1600 0 0 0 Mpp1
flabel comment s 4311 4824 4311 4824 0 FreeSans 1600 0 0 0 Mpp0
flabel comment s 2653 4824 2653 4824 0 FreeSans 1600 0 0 0 Mpp0
flabel comment s 995 4824 995 4824 0 FreeSans 1600 0 0 0 dum
flabel comment s 995 5324 995 5324 0 FreeSans 1600 0 0 0 dum
flabel comment s 2653 5324 2653 5324 0 FreeSans 1600 0 0 0 Mh0
flabel comment s 4311 5324 4311 5324 0 FreeSans 1600 0 0 0 Mh0
flabel comment s 5969 5324 5969 5324 0 FreeSans 1600 0 0 0 Mh1
flabel comment s 7627 5324 7627 5324 0 FreeSans 1600 0 0 0 Mh1
flabel comment s 9285 5324 9285 5324 0 FreeSans 1600 0 0 0 dum
flabel comment s 9285 7324 9285 7324 0 FreeSans 1600 0 0 0 dum
flabel comment s 7627 7324 7627 7324 0 FreeSans 1600 0 0 0 Mld0
flabel comment s 5969 7324 5969 7324 0 FreeSans 1600 0 0 0 Mld0
flabel comment s 4311 7324 4311 7324 0 FreeSans 1600 0 0 0 Mld1
flabel comment s 2653 7324 2653 7324 0 FreeSans 1600 0 0 0 Mld1
flabel comment s 995 7324 995 7324 0 FreeSans 1600 0 0 0 dum
flabel comment s -452 6161 -452 6161 0 FreeSans 800 0 0 0 Mt0
flabel comment s -452 6526 -452 6526 0 FreeSans 800 0 0 0 Minv1
flabel comment s -452 6891 -452 6891 0 FreeSans 800 0 0 0 Ml3
flabel comment s -452 7256 -452 7256 0 FreeSans 800 0 0 0 Ml4
flabel comment s -479 3464 -479 3464 0 FreeSans 800 0 0 0 Ml2
flabel comment s -479 4559 -479 4559 0 FreeSans 800 0 0 0 Minv0
flabel comment s -479 4924 -479 4924 0 FreeSans 800 0 0 0 Mt1
flabel comment s -488 4217 -488 4217 0 FreeSans 800 0 0 0 Ml0
flabel comment s -488 3861 -488 3861 0 FreeSans 800 0 0 0 Ml1
flabel metal3 -624 5359 -624 5359 7 FreeSans 1200 0 0 0 ibias
port 2 w
flabel metal2 -765 5650 -765 5650 7 FreeSans 1200 0 0 0 ena
port 4 w
flabel metal2 -205 5718 -205 5718 7 FreeSans 800 0 0 0 ena_b
flabel metal2 6740 4230 6740 4230 7 FreeSans 800 0 0 0 n0
flabel metal3 1755 2317 1755 2317 7 FreeSans 800 0 0 0 vnn
flabel metal3 1766 2517 1766 2517 7 FreeSans 800 0 0 0 vt
flabel metal3 1766 2717 1766 2717 7 FreeSans 800 0 0 0 vpp
flabel metal3 1766 2917 1766 2917 7 FreeSans 1200 0 0 0 vinn
port 5 w
flabel metal3 1766 3117 1766 3117 7 FreeSans 1200 0 0 0 vinp
port 6 w
flabel metal3 -619 7860 -619 7860 7 FreeSans 1200 0 0 0 avdd
port 1 w
flabel metal3 97 -77 97 -77 7 FreeSans 1200 0 0 0 avss
port 7 w
flabel metal2 10704 3729 10704 3729 3 FreeSans 800 0 0 0 n1
flabel metal3 10472 6132 10472 6132 1 FreeSans 1200 0 0 0 out
port 3 n
<< end >>
