magic
tech sky130A
magscale 1 2
timestamp 1711568248
<< nwell >>
rect -6861 -339 6861 339
<< mvpmos >>
rect -6603 -42 -5003 42
rect -4945 -42 -3345 42
rect -3287 -42 -1687 42
rect -1629 -42 -29 42
rect 29 -42 1629 42
rect 1687 -42 3287 42
rect 3345 -42 4945 42
rect 5003 -42 6603 42
<< mvpdiff >>
rect -6661 30 -6603 42
rect -6661 -30 -6649 30
rect -6615 -30 -6603 30
rect -6661 -42 -6603 -30
rect -5003 30 -4945 42
rect -5003 -30 -4991 30
rect -4957 -30 -4945 30
rect -5003 -42 -4945 -30
rect -3345 30 -3287 42
rect -3345 -30 -3333 30
rect -3299 -30 -3287 30
rect -3345 -42 -3287 -30
rect -1687 30 -1629 42
rect -1687 -30 -1675 30
rect -1641 -30 -1629 30
rect -1687 -42 -1629 -30
rect -29 30 29 42
rect -29 -30 -17 30
rect 17 -30 29 30
rect -29 -42 29 -30
rect 1629 30 1687 42
rect 1629 -30 1641 30
rect 1675 -30 1687 30
rect 1629 -42 1687 -30
rect 3287 30 3345 42
rect 3287 -30 3299 30
rect 3333 -30 3345 30
rect 3287 -42 3345 -30
rect 4945 30 5003 42
rect 4945 -30 4957 30
rect 4991 -30 5003 30
rect 4945 -42 5003 -30
rect 6603 30 6661 42
rect 6603 -30 6615 30
rect 6649 -30 6661 30
rect 6603 -42 6661 -30
<< mvpdiffc >>
rect -6649 -30 -6615 30
rect -4991 -30 -4957 30
rect -3333 -30 -3299 30
rect -1675 -30 -1641 30
rect -17 -30 17 30
rect 1641 -30 1675 30
rect 3299 -30 3333 30
rect 4957 -30 4991 30
rect 6615 -30 6649 30
<< mvnsubdiff >>
rect -6795 261 6795 273
rect -6795 227 -6687 261
rect 6687 227 6795 261
rect -6795 215 6795 227
rect -6795 165 -6737 215
rect -6795 -165 -6783 165
rect -6749 -165 -6737 165
rect 6737 165 6795 215
rect -6795 -215 -6737 -165
rect 6737 -165 6749 165
rect 6783 -165 6795 165
rect 6737 -215 6795 -165
rect -6795 -227 6795 -215
rect -6795 -261 -6687 -227
rect 6687 -261 6795 -227
rect -6795 -273 6795 -261
<< mvnsubdiffcont >>
rect -6687 227 6687 261
rect -6783 -165 -6749 165
rect 6749 -165 6783 165
rect -6687 -261 6687 -227
<< poly >>
rect -6603 123 -5003 139
rect -6603 89 -6587 123
rect -5019 89 -5003 123
rect -6603 42 -5003 89
rect -4945 123 -3345 139
rect -4945 89 -4929 123
rect -3361 89 -3345 123
rect -4945 42 -3345 89
rect -3287 123 -1687 139
rect -3287 89 -3271 123
rect -1703 89 -1687 123
rect -3287 42 -1687 89
rect -1629 123 -29 139
rect -1629 89 -1613 123
rect -45 89 -29 123
rect -1629 42 -29 89
rect 29 123 1629 139
rect 29 89 45 123
rect 1613 89 1629 123
rect 29 42 1629 89
rect 1687 123 3287 139
rect 1687 89 1703 123
rect 3271 89 3287 123
rect 1687 42 3287 89
rect 3345 123 4945 139
rect 3345 89 3361 123
rect 4929 89 4945 123
rect 3345 42 4945 89
rect 5003 123 6603 139
rect 5003 89 5019 123
rect 6587 89 6603 123
rect 5003 42 6603 89
rect -6603 -89 -5003 -42
rect -6603 -123 -6587 -89
rect -5019 -123 -5003 -89
rect -6603 -139 -5003 -123
rect -4945 -89 -3345 -42
rect -4945 -123 -4929 -89
rect -3361 -123 -3345 -89
rect -4945 -139 -3345 -123
rect -3287 -89 -1687 -42
rect -3287 -123 -3271 -89
rect -1703 -123 -1687 -89
rect -3287 -139 -1687 -123
rect -1629 -89 -29 -42
rect -1629 -123 -1613 -89
rect -45 -123 -29 -89
rect -1629 -139 -29 -123
rect 29 -89 1629 -42
rect 29 -123 45 -89
rect 1613 -123 1629 -89
rect 29 -139 1629 -123
rect 1687 -89 3287 -42
rect 1687 -123 1703 -89
rect 3271 -123 3287 -89
rect 1687 -139 3287 -123
rect 3345 -89 4945 -42
rect 3345 -123 3361 -89
rect 4929 -123 4945 -89
rect 3345 -139 4945 -123
rect 5003 -89 6603 -42
rect 5003 -123 5019 -89
rect 6587 -123 6603 -89
rect 5003 -139 6603 -123
<< polycont >>
rect -6587 89 -5019 123
rect -4929 89 -3361 123
rect -3271 89 -1703 123
rect -1613 89 -45 123
rect 45 89 1613 123
rect 1703 89 3271 123
rect 3361 89 4929 123
rect 5019 89 6587 123
rect -6587 -123 -5019 -89
rect -4929 -123 -3361 -89
rect -3271 -123 -1703 -89
rect -1613 -123 -45 -89
rect 45 -123 1613 -89
rect 1703 -123 3271 -89
rect 3361 -123 4929 -89
rect 5019 -123 6587 -89
<< locali >>
rect -6783 227 -6687 261
rect 6687 227 6783 261
rect -6783 165 -6749 227
rect 6749 165 6783 227
rect -6603 89 -6587 123
rect -5019 89 -5003 123
rect -4945 89 -4929 123
rect -3361 89 -3345 123
rect -3287 89 -3271 123
rect -1703 89 -1687 123
rect -1629 89 -1613 123
rect -45 89 -29 123
rect 29 89 45 123
rect 1613 89 1629 123
rect 1687 89 1703 123
rect 3271 89 3287 123
rect 3345 89 3361 123
rect 4929 89 4945 123
rect 5003 89 5019 123
rect 6587 89 6603 123
rect -6649 30 -6615 46
rect -6649 -46 -6615 -30
rect -4991 30 -4957 46
rect -4991 -46 -4957 -30
rect -3333 30 -3299 46
rect -3333 -46 -3299 -30
rect -1675 30 -1641 46
rect -1675 -46 -1641 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 1641 30 1675 46
rect 1641 -46 1675 -30
rect 3299 30 3333 46
rect 3299 -46 3333 -30
rect 4957 30 4991 46
rect 4957 -46 4991 -30
rect 6615 30 6649 46
rect 6615 -46 6649 -30
rect -6603 -123 -6587 -89
rect -5019 -123 -5003 -89
rect -4945 -123 -4929 -89
rect -3361 -123 -3345 -89
rect -3287 -123 -3271 -89
rect -1703 -123 -1687 -89
rect -1629 -123 -1613 -89
rect -45 -123 -29 -89
rect 29 -123 45 -89
rect 1613 -123 1629 -89
rect 1687 -123 1703 -89
rect 3271 -123 3287 -89
rect 3345 -123 3361 -89
rect 4929 -123 4945 -89
rect 5003 -123 5019 -89
rect 6587 -123 6603 -89
rect -6783 -227 -6749 -165
rect 6749 -227 6783 -165
rect -6783 -261 -6687 -227
rect 6687 -261 6783 -227
<< viali >>
rect -6587 89 -5019 123
rect -4929 89 -3361 123
rect -3271 89 -1703 123
rect -1613 89 -45 123
rect 45 89 1613 123
rect 1703 89 3271 123
rect 3361 89 4929 123
rect 5019 89 6587 123
rect -6649 -30 -6615 30
rect -4991 -30 -4957 30
rect -3333 -30 -3299 30
rect -1675 -30 -1641 30
rect -17 -30 17 30
rect 1641 -30 1675 30
rect 3299 -30 3333 30
rect 4957 -30 4991 30
rect 6615 -30 6649 30
rect -6587 -123 -5019 -89
rect -4929 -123 -3361 -89
rect -3271 -123 -1703 -89
rect -1613 -123 -45 -89
rect 45 -123 1613 -89
rect 1703 -123 3271 -89
rect 3361 -123 4929 -89
rect 5019 -123 6587 -89
<< metal1 >>
rect -6599 123 -5007 129
rect -6599 89 -6587 123
rect -5019 89 -5007 123
rect -6599 83 -5007 89
rect -4941 123 -3349 129
rect -4941 89 -4929 123
rect -3361 89 -3349 123
rect -4941 83 -3349 89
rect -3283 123 -1691 129
rect -3283 89 -3271 123
rect -1703 89 -1691 123
rect -3283 83 -1691 89
rect -1625 123 -33 129
rect -1625 89 -1613 123
rect -45 89 -33 123
rect -1625 83 -33 89
rect 33 123 1625 129
rect 33 89 45 123
rect 1613 89 1625 123
rect 33 83 1625 89
rect 1691 123 3283 129
rect 1691 89 1703 123
rect 3271 89 3283 123
rect 1691 83 3283 89
rect 3349 123 4941 129
rect 3349 89 3361 123
rect 4929 89 4941 123
rect 3349 83 4941 89
rect 5007 123 6599 129
rect 5007 89 5019 123
rect 6587 89 6599 123
rect 5007 83 6599 89
rect -6655 30 -6609 42
rect -6655 -30 -6649 30
rect -6615 -30 -6609 30
rect -6655 -42 -6609 -30
rect -4997 30 -4951 42
rect -4997 -30 -4991 30
rect -4957 -30 -4951 30
rect -4997 -42 -4951 -30
rect -3339 30 -3293 42
rect -3339 -30 -3333 30
rect -3299 -30 -3293 30
rect -3339 -42 -3293 -30
rect -1681 30 -1635 42
rect -1681 -30 -1675 30
rect -1641 -30 -1635 30
rect -1681 -42 -1635 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 1635 30 1681 42
rect 1635 -30 1641 30
rect 1675 -30 1681 30
rect 1635 -42 1681 -30
rect 3293 30 3339 42
rect 3293 -30 3299 30
rect 3333 -30 3339 30
rect 3293 -42 3339 -30
rect 4951 30 4997 42
rect 4951 -30 4957 30
rect 4991 -30 4997 30
rect 4951 -42 4997 -30
rect 6609 30 6655 42
rect 6609 -30 6615 30
rect 6649 -30 6655 30
rect 6609 -42 6655 -30
rect -6599 -89 -5007 -83
rect -6599 -123 -6587 -89
rect -5019 -123 -5007 -89
rect -6599 -129 -5007 -123
rect -4941 -89 -3349 -83
rect -4941 -123 -4929 -89
rect -3361 -123 -3349 -89
rect -4941 -129 -3349 -123
rect -3283 -89 -1691 -83
rect -3283 -123 -3271 -89
rect -1703 -123 -1691 -89
rect -3283 -129 -1691 -123
rect -1625 -89 -33 -83
rect -1625 -123 -1613 -89
rect -45 -123 -33 -89
rect -1625 -129 -33 -123
rect 33 -89 1625 -83
rect 33 -123 45 -89
rect 1613 -123 1625 -89
rect 33 -129 1625 -123
rect 1691 -89 3283 -83
rect 1691 -123 1703 -89
rect 3271 -123 3283 -89
rect 1691 -129 3283 -123
rect 3349 -89 4941 -83
rect 3349 -123 3361 -89
rect 4929 -123 4941 -89
rect 3349 -129 4941 -123
rect 5007 -89 6599 -83
rect 5007 -123 5019 -89
rect 6587 -123 6599 -89
rect 5007 -129 6599 -123
<< properties >>
string FIXED_BBOX -6766 -244 6766 244
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 8.0 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
