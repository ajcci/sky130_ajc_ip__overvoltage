magic
tech sky130A
magscale 1 2
timestamp 1712105914
<< pwell >>
rect -5173 -1976 5173 1976
<< mvnmos >>
rect -4945 718 -3345 1718
rect -3287 718 -1687 1718
rect -1629 718 -29 1718
rect 29 718 1629 1718
rect 1687 718 3287 1718
rect 3345 718 4945 1718
rect -4945 -500 -3345 500
rect -3287 -500 -1687 500
rect -1629 -500 -29 500
rect 29 -500 1629 500
rect 1687 -500 3287 500
rect 3345 -500 4945 500
rect -4945 -1718 -3345 -718
rect -3287 -1718 -1687 -718
rect -1629 -1718 -29 -718
rect 29 -1718 1629 -718
rect 1687 -1718 3287 -718
rect 3345 -1718 4945 -718
<< mvndiff >>
rect -5003 1706 -4945 1718
rect -5003 730 -4991 1706
rect -4957 730 -4945 1706
rect -5003 718 -4945 730
rect -3345 1706 -3287 1718
rect -3345 730 -3333 1706
rect -3299 730 -3287 1706
rect -3345 718 -3287 730
rect -1687 1706 -1629 1718
rect -1687 730 -1675 1706
rect -1641 730 -1629 1706
rect -1687 718 -1629 730
rect -29 1706 29 1718
rect -29 730 -17 1706
rect 17 730 29 1706
rect -29 718 29 730
rect 1629 1706 1687 1718
rect 1629 730 1641 1706
rect 1675 730 1687 1706
rect 1629 718 1687 730
rect 3287 1706 3345 1718
rect 3287 730 3299 1706
rect 3333 730 3345 1706
rect 3287 718 3345 730
rect 4945 1706 5003 1718
rect 4945 730 4957 1706
rect 4991 730 5003 1706
rect 4945 718 5003 730
rect -5003 488 -4945 500
rect -5003 -488 -4991 488
rect -4957 -488 -4945 488
rect -5003 -500 -4945 -488
rect -3345 488 -3287 500
rect -3345 -488 -3333 488
rect -3299 -488 -3287 488
rect -3345 -500 -3287 -488
rect -1687 488 -1629 500
rect -1687 -488 -1675 488
rect -1641 -488 -1629 488
rect -1687 -500 -1629 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 1629 488 1687 500
rect 1629 -488 1641 488
rect 1675 -488 1687 488
rect 1629 -500 1687 -488
rect 3287 488 3345 500
rect 3287 -488 3299 488
rect 3333 -488 3345 488
rect 3287 -500 3345 -488
rect 4945 488 5003 500
rect 4945 -488 4957 488
rect 4991 -488 5003 488
rect 4945 -500 5003 -488
rect -5003 -730 -4945 -718
rect -5003 -1706 -4991 -730
rect -4957 -1706 -4945 -730
rect -5003 -1718 -4945 -1706
rect -3345 -730 -3287 -718
rect -3345 -1706 -3333 -730
rect -3299 -1706 -3287 -730
rect -3345 -1718 -3287 -1706
rect -1687 -730 -1629 -718
rect -1687 -1706 -1675 -730
rect -1641 -1706 -1629 -730
rect -1687 -1718 -1629 -1706
rect -29 -730 29 -718
rect -29 -1706 -17 -730
rect 17 -1706 29 -730
rect -29 -1718 29 -1706
rect 1629 -730 1687 -718
rect 1629 -1706 1641 -730
rect 1675 -1706 1687 -730
rect 1629 -1718 1687 -1706
rect 3287 -730 3345 -718
rect 3287 -1706 3299 -730
rect 3333 -1706 3345 -730
rect 3287 -1718 3345 -1706
rect 4945 -730 5003 -718
rect 4945 -1706 4957 -730
rect 4991 -1706 5003 -730
rect 4945 -1718 5003 -1706
<< mvndiffc >>
rect -4991 730 -4957 1706
rect -3333 730 -3299 1706
rect -1675 730 -1641 1706
rect -17 730 17 1706
rect 1641 730 1675 1706
rect 3299 730 3333 1706
rect 4957 730 4991 1706
rect -4991 -488 -4957 488
rect -3333 -488 -3299 488
rect -1675 -488 -1641 488
rect -17 -488 17 488
rect 1641 -488 1675 488
rect 3299 -488 3333 488
rect 4957 -488 4991 488
rect -4991 -1706 -4957 -730
rect -3333 -1706 -3299 -730
rect -1675 -1706 -1641 -730
rect -17 -1706 17 -730
rect 1641 -1706 1675 -730
rect 3299 -1706 3333 -730
rect 4957 -1706 4991 -730
<< mvpsubdiff >>
rect -5137 1928 5137 1940
rect -5137 1894 -5029 1928
rect 5029 1894 5137 1928
rect -5137 1882 5137 1894
rect -5137 1832 -5079 1882
rect -5137 -1832 -5125 1832
rect -5091 -1832 -5079 1832
rect 5079 1832 5137 1882
rect -5137 -1882 -5079 -1832
rect 5079 -1832 5091 1832
rect 5125 -1832 5137 1832
rect 5079 -1882 5137 -1832
rect -5137 -1894 5137 -1882
rect -5137 -1928 -5029 -1894
rect 5029 -1928 5137 -1894
rect -5137 -1940 5137 -1928
<< mvpsubdiffcont >>
rect -5029 1894 5029 1928
rect -5125 -1832 -5091 1832
rect 5091 -1832 5125 1832
rect -5029 -1928 5029 -1894
<< poly >>
rect -4945 1790 -3345 1806
rect -4945 1756 -4929 1790
rect -3361 1756 -3345 1790
rect -4945 1718 -3345 1756
rect -3287 1790 -1687 1806
rect -3287 1756 -3271 1790
rect -1703 1756 -1687 1790
rect -3287 1718 -1687 1756
rect -1629 1790 -29 1806
rect -1629 1756 -1613 1790
rect -45 1756 -29 1790
rect -1629 1718 -29 1756
rect 29 1790 1629 1806
rect 29 1756 45 1790
rect 1613 1756 1629 1790
rect 29 1718 1629 1756
rect 1687 1790 3287 1806
rect 1687 1756 1703 1790
rect 3271 1756 3287 1790
rect 1687 1718 3287 1756
rect 3345 1790 4945 1806
rect 3345 1756 3361 1790
rect 4929 1756 4945 1790
rect 3345 1718 4945 1756
rect -4945 680 -3345 718
rect -4945 646 -4929 680
rect -3361 646 -3345 680
rect -4945 630 -3345 646
rect -3287 680 -1687 718
rect -3287 646 -3271 680
rect -1703 646 -1687 680
rect -3287 630 -1687 646
rect -1629 680 -29 718
rect -1629 646 -1613 680
rect -45 646 -29 680
rect -1629 630 -29 646
rect 29 680 1629 718
rect 29 646 45 680
rect 1613 646 1629 680
rect 29 630 1629 646
rect 1687 680 3287 718
rect 1687 646 1703 680
rect 3271 646 3287 680
rect 1687 630 3287 646
rect 3345 680 4945 718
rect 3345 646 3361 680
rect 4929 646 4945 680
rect 3345 630 4945 646
rect -4945 572 -3345 588
rect -4945 538 -4929 572
rect -3361 538 -3345 572
rect -4945 500 -3345 538
rect -3287 572 -1687 588
rect -3287 538 -3271 572
rect -1703 538 -1687 572
rect -3287 500 -1687 538
rect -1629 572 -29 588
rect -1629 538 -1613 572
rect -45 538 -29 572
rect -1629 500 -29 538
rect 29 572 1629 588
rect 29 538 45 572
rect 1613 538 1629 572
rect 29 500 1629 538
rect 1687 572 3287 588
rect 1687 538 1703 572
rect 3271 538 3287 572
rect 1687 500 3287 538
rect 3345 572 4945 588
rect 3345 538 3361 572
rect 4929 538 4945 572
rect 3345 500 4945 538
rect -4945 -538 -3345 -500
rect -4945 -572 -4929 -538
rect -3361 -572 -3345 -538
rect -4945 -588 -3345 -572
rect -3287 -538 -1687 -500
rect -3287 -572 -3271 -538
rect -1703 -572 -1687 -538
rect -3287 -588 -1687 -572
rect -1629 -538 -29 -500
rect -1629 -572 -1613 -538
rect -45 -572 -29 -538
rect -1629 -588 -29 -572
rect 29 -538 1629 -500
rect 29 -572 45 -538
rect 1613 -572 1629 -538
rect 29 -588 1629 -572
rect 1687 -538 3287 -500
rect 1687 -572 1703 -538
rect 3271 -572 3287 -538
rect 1687 -588 3287 -572
rect 3345 -538 4945 -500
rect 3345 -572 3361 -538
rect 4929 -572 4945 -538
rect 3345 -588 4945 -572
rect -4945 -646 -3345 -630
rect -4945 -680 -4929 -646
rect -3361 -680 -3345 -646
rect -4945 -718 -3345 -680
rect -3287 -646 -1687 -630
rect -3287 -680 -3271 -646
rect -1703 -680 -1687 -646
rect -3287 -718 -1687 -680
rect -1629 -646 -29 -630
rect -1629 -680 -1613 -646
rect -45 -680 -29 -646
rect -1629 -718 -29 -680
rect 29 -646 1629 -630
rect 29 -680 45 -646
rect 1613 -680 1629 -646
rect 29 -718 1629 -680
rect 1687 -646 3287 -630
rect 1687 -680 1703 -646
rect 3271 -680 3287 -646
rect 1687 -718 3287 -680
rect 3345 -646 4945 -630
rect 3345 -680 3361 -646
rect 4929 -680 4945 -646
rect 3345 -718 4945 -680
rect -4945 -1756 -3345 -1718
rect -4945 -1790 -4929 -1756
rect -3361 -1790 -3345 -1756
rect -4945 -1806 -3345 -1790
rect -3287 -1756 -1687 -1718
rect -3287 -1790 -3271 -1756
rect -1703 -1790 -1687 -1756
rect -3287 -1806 -1687 -1790
rect -1629 -1756 -29 -1718
rect -1629 -1790 -1613 -1756
rect -45 -1790 -29 -1756
rect -1629 -1806 -29 -1790
rect 29 -1756 1629 -1718
rect 29 -1790 45 -1756
rect 1613 -1790 1629 -1756
rect 29 -1806 1629 -1790
rect 1687 -1756 3287 -1718
rect 1687 -1790 1703 -1756
rect 3271 -1790 3287 -1756
rect 1687 -1806 3287 -1790
rect 3345 -1756 4945 -1718
rect 3345 -1790 3361 -1756
rect 4929 -1790 4945 -1756
rect 3345 -1806 4945 -1790
<< polycont >>
rect -4929 1756 -3361 1790
rect -3271 1756 -1703 1790
rect -1613 1756 -45 1790
rect 45 1756 1613 1790
rect 1703 1756 3271 1790
rect 3361 1756 4929 1790
rect -4929 646 -3361 680
rect -3271 646 -1703 680
rect -1613 646 -45 680
rect 45 646 1613 680
rect 1703 646 3271 680
rect 3361 646 4929 680
rect -4929 538 -3361 572
rect -3271 538 -1703 572
rect -1613 538 -45 572
rect 45 538 1613 572
rect 1703 538 3271 572
rect 3361 538 4929 572
rect -4929 -572 -3361 -538
rect -3271 -572 -1703 -538
rect -1613 -572 -45 -538
rect 45 -572 1613 -538
rect 1703 -572 3271 -538
rect 3361 -572 4929 -538
rect -4929 -680 -3361 -646
rect -3271 -680 -1703 -646
rect -1613 -680 -45 -646
rect 45 -680 1613 -646
rect 1703 -680 3271 -646
rect 3361 -680 4929 -646
rect -4929 -1790 -3361 -1756
rect -3271 -1790 -1703 -1756
rect -1613 -1790 -45 -1756
rect 45 -1790 1613 -1756
rect 1703 -1790 3271 -1756
rect 3361 -1790 4929 -1756
<< locali >>
rect -5125 1894 -5029 1928
rect 5029 1894 5125 1928
rect -5125 1832 -5091 1894
rect 5091 1832 5125 1894
rect -4945 1756 -4929 1790
rect -3361 1756 -3345 1790
rect -3287 1756 -3271 1790
rect -1703 1756 -1687 1790
rect -1629 1756 -1613 1790
rect -45 1756 -29 1790
rect 29 1756 45 1790
rect 1613 1756 1629 1790
rect 1687 1756 1703 1790
rect 3271 1756 3287 1790
rect 3345 1756 3361 1790
rect 4929 1756 4945 1790
rect -4991 1706 -4957 1722
rect -4991 714 -4957 730
rect -3333 1706 -3299 1722
rect -3333 714 -3299 730
rect -1675 1706 -1641 1722
rect -1675 714 -1641 730
rect -17 1706 17 1722
rect -17 714 17 730
rect 1641 1706 1675 1722
rect 1641 714 1675 730
rect 3299 1706 3333 1722
rect 3299 714 3333 730
rect 4957 1706 4991 1722
rect 4957 714 4991 730
rect -4945 646 -4929 680
rect -3361 646 -3345 680
rect -3287 646 -3271 680
rect -1703 646 -1687 680
rect -1629 646 -1613 680
rect -45 646 -29 680
rect 29 646 45 680
rect 1613 646 1629 680
rect 1687 646 1703 680
rect 3271 646 3287 680
rect 3345 646 3361 680
rect 4929 646 4945 680
rect -4945 538 -4929 572
rect -3361 538 -3345 572
rect -3287 538 -3271 572
rect -1703 538 -1687 572
rect -1629 538 -1613 572
rect -45 538 -29 572
rect 29 538 45 572
rect 1613 538 1629 572
rect 1687 538 1703 572
rect 3271 538 3287 572
rect 3345 538 3361 572
rect 4929 538 4945 572
rect -4991 488 -4957 504
rect -4991 -504 -4957 -488
rect -3333 488 -3299 504
rect -3333 -504 -3299 -488
rect -1675 488 -1641 504
rect -1675 -504 -1641 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 1641 488 1675 504
rect 1641 -504 1675 -488
rect 3299 488 3333 504
rect 3299 -504 3333 -488
rect 4957 488 4991 504
rect 4957 -504 4991 -488
rect -4945 -572 -4929 -538
rect -3361 -572 -3345 -538
rect -3287 -572 -3271 -538
rect -1703 -572 -1687 -538
rect -1629 -572 -1613 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 1613 -572 1629 -538
rect 1687 -572 1703 -538
rect 3271 -572 3287 -538
rect 3345 -572 3361 -538
rect 4929 -572 4945 -538
rect -4945 -680 -4929 -646
rect -3361 -680 -3345 -646
rect -3287 -680 -3271 -646
rect -1703 -680 -1687 -646
rect -1629 -680 -1613 -646
rect -45 -680 -29 -646
rect 29 -680 45 -646
rect 1613 -680 1629 -646
rect 1687 -680 1703 -646
rect 3271 -680 3287 -646
rect 3345 -680 3361 -646
rect 4929 -680 4945 -646
rect -4991 -730 -4957 -714
rect -4991 -1722 -4957 -1706
rect -3333 -730 -3299 -714
rect -3333 -1722 -3299 -1706
rect -1675 -730 -1641 -714
rect -1675 -1722 -1641 -1706
rect -17 -730 17 -714
rect -17 -1722 17 -1706
rect 1641 -730 1675 -714
rect 1641 -1722 1675 -1706
rect 3299 -730 3333 -714
rect 3299 -1722 3333 -1706
rect 4957 -730 4991 -714
rect 4957 -1722 4991 -1706
rect -4945 -1790 -4929 -1756
rect -3361 -1790 -3345 -1756
rect -3287 -1790 -3271 -1756
rect -1703 -1790 -1687 -1756
rect -1629 -1790 -1613 -1756
rect -45 -1790 -29 -1756
rect 29 -1790 45 -1756
rect 1613 -1790 1629 -1756
rect 1687 -1790 1703 -1756
rect 3271 -1790 3287 -1756
rect 3345 -1790 3361 -1756
rect 4929 -1790 4945 -1756
rect -5125 -1894 -5091 -1832
rect 5091 -1894 5125 -1832
rect -5125 -1928 -5029 -1894
rect 5029 -1928 5125 -1894
<< viali >>
rect -4929 1756 -3361 1790
rect -3271 1756 -1703 1790
rect -1613 1756 -45 1790
rect 45 1756 1613 1790
rect 1703 1756 3271 1790
rect 3361 1756 4929 1790
rect -4991 730 -4957 1706
rect -3333 730 -3299 1706
rect -1675 730 -1641 1706
rect -17 730 17 1706
rect 1641 730 1675 1706
rect 3299 730 3333 1706
rect 4957 730 4991 1706
rect -4929 646 -3361 680
rect -3271 646 -1703 680
rect -1613 646 -45 680
rect 45 646 1613 680
rect 1703 646 3271 680
rect 3361 646 4929 680
rect -4929 538 -3361 572
rect -3271 538 -1703 572
rect -1613 538 -45 572
rect 45 538 1613 572
rect 1703 538 3271 572
rect 3361 538 4929 572
rect -4991 -488 -4957 488
rect -3333 -488 -3299 488
rect -1675 -488 -1641 488
rect -17 -488 17 488
rect 1641 -488 1675 488
rect 3299 -488 3333 488
rect 4957 -488 4991 488
rect -4929 -572 -3361 -538
rect -3271 -572 -1703 -538
rect -1613 -572 -45 -538
rect 45 -572 1613 -538
rect 1703 -572 3271 -538
rect 3361 -572 4929 -538
rect -4929 -680 -3361 -646
rect -3271 -680 -1703 -646
rect -1613 -680 -45 -646
rect 45 -680 1613 -646
rect 1703 -680 3271 -646
rect 3361 -680 4929 -646
rect -4991 -1706 -4957 -730
rect -3333 -1706 -3299 -730
rect -1675 -1706 -1641 -730
rect -17 -1706 17 -730
rect 1641 -1706 1675 -730
rect 3299 -1706 3333 -730
rect 4957 -1706 4991 -730
rect -4929 -1790 -3361 -1756
rect -3271 -1790 -1703 -1756
rect -1613 -1790 -45 -1756
rect 45 -1790 1613 -1756
rect 1703 -1790 3271 -1756
rect 3361 -1790 4929 -1756
<< metal1 >>
rect -4941 1790 -3349 1796
rect -4941 1756 -4929 1790
rect -3361 1756 -3349 1790
rect -4941 1750 -3349 1756
rect -3283 1790 -1691 1796
rect -3283 1756 -3271 1790
rect -1703 1756 -1691 1790
rect -3283 1750 -1691 1756
rect -1625 1790 -33 1796
rect -1625 1756 -1613 1790
rect -45 1756 -33 1790
rect -1625 1750 -33 1756
rect 33 1790 1625 1796
rect 33 1756 45 1790
rect 1613 1756 1625 1790
rect 33 1750 1625 1756
rect 1691 1790 3283 1796
rect 1691 1756 1703 1790
rect 3271 1756 3283 1790
rect 1691 1750 3283 1756
rect 3349 1790 4941 1796
rect 3349 1756 3361 1790
rect 4929 1756 4941 1790
rect 3349 1750 4941 1756
rect -4997 1706 -4951 1718
rect -4997 730 -4991 1706
rect -4957 730 -4951 1706
rect -4997 718 -4951 730
rect -3339 1706 -3293 1718
rect -3339 730 -3333 1706
rect -3299 730 -3293 1706
rect -3339 718 -3293 730
rect -1681 1706 -1635 1718
rect -1681 730 -1675 1706
rect -1641 730 -1635 1706
rect -1681 718 -1635 730
rect -23 1706 23 1718
rect -23 730 -17 1706
rect 17 730 23 1706
rect -23 718 23 730
rect 1635 1706 1681 1718
rect 1635 730 1641 1706
rect 1675 730 1681 1706
rect 1635 718 1681 730
rect 3293 1706 3339 1718
rect 3293 730 3299 1706
rect 3333 730 3339 1706
rect 3293 718 3339 730
rect 4951 1706 4997 1718
rect 4951 730 4957 1706
rect 4991 730 4997 1706
rect 4951 718 4997 730
rect -4941 680 -3349 686
rect -4941 646 -4929 680
rect -3361 646 -3349 680
rect -4941 640 -3349 646
rect -3283 680 -1691 686
rect -3283 646 -3271 680
rect -1703 646 -1691 680
rect -3283 640 -1691 646
rect -1625 680 -33 686
rect -1625 646 -1613 680
rect -45 646 -33 680
rect -1625 640 -33 646
rect 33 680 1625 686
rect 33 646 45 680
rect 1613 646 1625 680
rect 33 640 1625 646
rect 1691 680 3283 686
rect 1691 646 1703 680
rect 3271 646 3283 680
rect 1691 640 3283 646
rect 3349 680 4941 686
rect 3349 646 3361 680
rect 4929 646 4941 680
rect 3349 640 4941 646
rect -4941 572 -3349 578
rect -4941 538 -4929 572
rect -3361 538 -3349 572
rect -4941 532 -3349 538
rect -3283 572 -1691 578
rect -3283 538 -3271 572
rect -1703 538 -1691 572
rect -3283 532 -1691 538
rect -1625 572 -33 578
rect -1625 538 -1613 572
rect -45 538 -33 572
rect -1625 532 -33 538
rect 33 572 1625 578
rect 33 538 45 572
rect 1613 538 1625 572
rect 33 532 1625 538
rect 1691 572 3283 578
rect 1691 538 1703 572
rect 3271 538 3283 572
rect 1691 532 3283 538
rect 3349 572 4941 578
rect 3349 538 3361 572
rect 4929 538 4941 572
rect 3349 532 4941 538
rect -4997 488 -4951 500
rect -4997 -488 -4991 488
rect -4957 -488 -4951 488
rect -4997 -500 -4951 -488
rect -3339 488 -3293 500
rect -3339 -488 -3333 488
rect -3299 -488 -3293 488
rect -3339 -500 -3293 -488
rect -1681 488 -1635 500
rect -1681 -488 -1675 488
rect -1641 -488 -1635 488
rect -1681 -500 -1635 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 1635 488 1681 500
rect 1635 -488 1641 488
rect 1675 -488 1681 488
rect 1635 -500 1681 -488
rect 3293 488 3339 500
rect 3293 -488 3299 488
rect 3333 -488 3339 488
rect 3293 -500 3339 -488
rect 4951 488 4997 500
rect 4951 -488 4957 488
rect 4991 -488 4997 488
rect 4951 -500 4997 -488
rect -4941 -538 -3349 -532
rect -4941 -572 -4929 -538
rect -3361 -572 -3349 -538
rect -4941 -578 -3349 -572
rect -3283 -538 -1691 -532
rect -3283 -572 -3271 -538
rect -1703 -572 -1691 -538
rect -3283 -578 -1691 -572
rect -1625 -538 -33 -532
rect -1625 -572 -1613 -538
rect -45 -572 -33 -538
rect -1625 -578 -33 -572
rect 33 -538 1625 -532
rect 33 -572 45 -538
rect 1613 -572 1625 -538
rect 33 -578 1625 -572
rect 1691 -538 3283 -532
rect 1691 -572 1703 -538
rect 3271 -572 3283 -538
rect 1691 -578 3283 -572
rect 3349 -538 4941 -532
rect 3349 -572 3361 -538
rect 4929 -572 4941 -538
rect 3349 -578 4941 -572
rect -4941 -646 -3349 -640
rect -4941 -680 -4929 -646
rect -3361 -680 -3349 -646
rect -4941 -686 -3349 -680
rect -3283 -646 -1691 -640
rect -3283 -680 -3271 -646
rect -1703 -680 -1691 -646
rect -3283 -686 -1691 -680
rect -1625 -646 -33 -640
rect -1625 -680 -1613 -646
rect -45 -680 -33 -646
rect -1625 -686 -33 -680
rect 33 -646 1625 -640
rect 33 -680 45 -646
rect 1613 -680 1625 -646
rect 33 -686 1625 -680
rect 1691 -646 3283 -640
rect 1691 -680 1703 -646
rect 3271 -680 3283 -646
rect 1691 -686 3283 -680
rect 3349 -646 4941 -640
rect 3349 -680 3361 -646
rect 4929 -680 4941 -646
rect 3349 -686 4941 -680
rect -4997 -730 -4951 -718
rect -4997 -1706 -4991 -730
rect -4957 -1706 -4951 -730
rect -4997 -1718 -4951 -1706
rect -3339 -730 -3293 -718
rect -3339 -1706 -3333 -730
rect -3299 -1706 -3293 -730
rect -3339 -1718 -3293 -1706
rect -1681 -730 -1635 -718
rect -1681 -1706 -1675 -730
rect -1641 -1706 -1635 -730
rect -1681 -1718 -1635 -1706
rect -23 -730 23 -718
rect -23 -1706 -17 -730
rect 17 -1706 23 -730
rect -23 -1718 23 -1706
rect 1635 -730 1681 -718
rect 1635 -1706 1641 -730
rect 1675 -1706 1681 -730
rect 1635 -1718 1681 -1706
rect 3293 -730 3339 -718
rect 3293 -1706 3299 -730
rect 3333 -1706 3339 -730
rect 3293 -1718 3339 -1706
rect 4951 -730 4997 -718
rect 4951 -1706 4957 -730
rect 4991 -1706 4997 -730
rect 4951 -1718 4997 -1706
rect -4941 -1756 -3349 -1750
rect -4941 -1790 -4929 -1756
rect -3361 -1790 -3349 -1756
rect -4941 -1796 -3349 -1790
rect -3283 -1756 -1691 -1750
rect -3283 -1790 -3271 -1756
rect -1703 -1790 -1691 -1756
rect -3283 -1796 -1691 -1790
rect -1625 -1756 -33 -1750
rect -1625 -1790 -1613 -1756
rect -45 -1790 -33 -1756
rect -1625 -1796 -33 -1790
rect 33 -1756 1625 -1750
rect 33 -1790 45 -1756
rect 1613 -1790 1625 -1756
rect 33 -1796 1625 -1790
rect 1691 -1756 3283 -1750
rect 1691 -1790 1703 -1756
rect 3271 -1790 3283 -1756
rect 1691 -1796 3283 -1790
rect 3349 -1756 4941 -1750
rect 3349 -1790 3361 -1756
rect 4929 -1790 4941 -1756
rect 3349 -1796 4941 -1790
<< properties >>
string FIXED_BBOX -5108 -1911 5108 1911
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 8 m 3 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
