magic
tech sky130A
magscale 1 2
timestamp 1711568248
<< pwell >>
rect -13463 -300 13463 300
<< mvnmos >>
rect -13235 -42 -11635 42
rect -11577 -42 -9977 42
rect -9919 -42 -8319 42
rect -8261 -42 -6661 42
rect -6603 -42 -5003 42
rect -4945 -42 -3345 42
rect -3287 -42 -1687 42
rect -1629 -42 -29 42
rect 29 -42 1629 42
rect 1687 -42 3287 42
rect 3345 -42 4945 42
rect 5003 -42 6603 42
rect 6661 -42 8261 42
rect 8319 -42 9919 42
rect 9977 -42 11577 42
rect 11635 -42 13235 42
<< mvndiff >>
rect -13293 30 -13235 42
rect -13293 -30 -13281 30
rect -13247 -30 -13235 30
rect -13293 -42 -13235 -30
rect -11635 30 -11577 42
rect -11635 -30 -11623 30
rect -11589 -30 -11577 30
rect -11635 -42 -11577 -30
rect -9977 30 -9919 42
rect -9977 -30 -9965 30
rect -9931 -30 -9919 30
rect -9977 -42 -9919 -30
rect -8319 30 -8261 42
rect -8319 -30 -8307 30
rect -8273 -30 -8261 30
rect -8319 -42 -8261 -30
rect -6661 30 -6603 42
rect -6661 -30 -6649 30
rect -6615 -30 -6603 30
rect -6661 -42 -6603 -30
rect -5003 30 -4945 42
rect -5003 -30 -4991 30
rect -4957 -30 -4945 30
rect -5003 -42 -4945 -30
rect -3345 30 -3287 42
rect -3345 -30 -3333 30
rect -3299 -30 -3287 30
rect -3345 -42 -3287 -30
rect -1687 30 -1629 42
rect -1687 -30 -1675 30
rect -1641 -30 -1629 30
rect -1687 -42 -1629 -30
rect -29 30 29 42
rect -29 -30 -17 30
rect 17 -30 29 30
rect -29 -42 29 -30
rect 1629 30 1687 42
rect 1629 -30 1641 30
rect 1675 -30 1687 30
rect 1629 -42 1687 -30
rect 3287 30 3345 42
rect 3287 -30 3299 30
rect 3333 -30 3345 30
rect 3287 -42 3345 -30
rect 4945 30 5003 42
rect 4945 -30 4957 30
rect 4991 -30 5003 30
rect 4945 -42 5003 -30
rect 6603 30 6661 42
rect 6603 -30 6615 30
rect 6649 -30 6661 30
rect 6603 -42 6661 -30
rect 8261 30 8319 42
rect 8261 -30 8273 30
rect 8307 -30 8319 30
rect 8261 -42 8319 -30
rect 9919 30 9977 42
rect 9919 -30 9931 30
rect 9965 -30 9977 30
rect 9919 -42 9977 -30
rect 11577 30 11635 42
rect 11577 -30 11589 30
rect 11623 -30 11635 30
rect 11577 -42 11635 -30
rect 13235 30 13293 42
rect 13235 -30 13247 30
rect 13281 -30 13293 30
rect 13235 -42 13293 -30
<< mvndiffc >>
rect -13281 -30 -13247 30
rect -11623 -30 -11589 30
rect -9965 -30 -9931 30
rect -8307 -30 -8273 30
rect -6649 -30 -6615 30
rect -4991 -30 -4957 30
rect -3333 -30 -3299 30
rect -1675 -30 -1641 30
rect -17 -30 17 30
rect 1641 -30 1675 30
rect 3299 -30 3333 30
rect 4957 -30 4991 30
rect 6615 -30 6649 30
rect 8273 -30 8307 30
rect 9931 -30 9965 30
rect 11589 -30 11623 30
rect 13247 -30 13281 30
<< mvpsubdiff >>
rect -13427 252 13427 264
rect -13427 218 -13319 252
rect 13319 218 13427 252
rect -13427 206 13427 218
rect -13427 156 -13369 206
rect -13427 -156 -13415 156
rect -13381 -156 -13369 156
rect 13369 156 13427 206
rect -13427 -206 -13369 -156
rect 13369 -156 13381 156
rect 13415 -156 13427 156
rect 13369 -206 13427 -156
rect -13427 -218 13427 -206
rect -13427 -252 -13319 -218
rect 13319 -252 13427 -218
rect -13427 -264 13427 -252
<< mvpsubdiffcont >>
rect -13319 218 13319 252
rect -13415 -156 -13381 156
rect 13381 -156 13415 156
rect -13319 -252 13319 -218
<< poly >>
rect -13235 114 -11635 130
rect -13235 80 -13219 114
rect -11651 80 -11635 114
rect -13235 42 -11635 80
rect -11577 114 -9977 130
rect -11577 80 -11561 114
rect -9993 80 -9977 114
rect -11577 42 -9977 80
rect -9919 114 -8319 130
rect -9919 80 -9903 114
rect -8335 80 -8319 114
rect -9919 42 -8319 80
rect -8261 114 -6661 130
rect -8261 80 -8245 114
rect -6677 80 -6661 114
rect -8261 42 -6661 80
rect -6603 114 -5003 130
rect -6603 80 -6587 114
rect -5019 80 -5003 114
rect -6603 42 -5003 80
rect -4945 114 -3345 130
rect -4945 80 -4929 114
rect -3361 80 -3345 114
rect -4945 42 -3345 80
rect -3287 114 -1687 130
rect -3287 80 -3271 114
rect -1703 80 -1687 114
rect -3287 42 -1687 80
rect -1629 114 -29 130
rect -1629 80 -1613 114
rect -45 80 -29 114
rect -1629 42 -29 80
rect 29 114 1629 130
rect 29 80 45 114
rect 1613 80 1629 114
rect 29 42 1629 80
rect 1687 114 3287 130
rect 1687 80 1703 114
rect 3271 80 3287 114
rect 1687 42 3287 80
rect 3345 114 4945 130
rect 3345 80 3361 114
rect 4929 80 4945 114
rect 3345 42 4945 80
rect 5003 114 6603 130
rect 5003 80 5019 114
rect 6587 80 6603 114
rect 5003 42 6603 80
rect 6661 114 8261 130
rect 6661 80 6677 114
rect 8245 80 8261 114
rect 6661 42 8261 80
rect 8319 114 9919 130
rect 8319 80 8335 114
rect 9903 80 9919 114
rect 8319 42 9919 80
rect 9977 114 11577 130
rect 9977 80 9993 114
rect 11561 80 11577 114
rect 9977 42 11577 80
rect 11635 114 13235 130
rect 11635 80 11651 114
rect 13219 80 13235 114
rect 11635 42 13235 80
rect -13235 -80 -11635 -42
rect -13235 -114 -13219 -80
rect -11651 -114 -11635 -80
rect -13235 -130 -11635 -114
rect -11577 -80 -9977 -42
rect -11577 -114 -11561 -80
rect -9993 -114 -9977 -80
rect -11577 -130 -9977 -114
rect -9919 -80 -8319 -42
rect -9919 -114 -9903 -80
rect -8335 -114 -8319 -80
rect -9919 -130 -8319 -114
rect -8261 -80 -6661 -42
rect -8261 -114 -8245 -80
rect -6677 -114 -6661 -80
rect -8261 -130 -6661 -114
rect -6603 -80 -5003 -42
rect -6603 -114 -6587 -80
rect -5019 -114 -5003 -80
rect -6603 -130 -5003 -114
rect -4945 -80 -3345 -42
rect -4945 -114 -4929 -80
rect -3361 -114 -3345 -80
rect -4945 -130 -3345 -114
rect -3287 -80 -1687 -42
rect -3287 -114 -3271 -80
rect -1703 -114 -1687 -80
rect -3287 -130 -1687 -114
rect -1629 -80 -29 -42
rect -1629 -114 -1613 -80
rect -45 -114 -29 -80
rect -1629 -130 -29 -114
rect 29 -80 1629 -42
rect 29 -114 45 -80
rect 1613 -114 1629 -80
rect 29 -130 1629 -114
rect 1687 -80 3287 -42
rect 1687 -114 1703 -80
rect 3271 -114 3287 -80
rect 1687 -130 3287 -114
rect 3345 -80 4945 -42
rect 3345 -114 3361 -80
rect 4929 -114 4945 -80
rect 3345 -130 4945 -114
rect 5003 -80 6603 -42
rect 5003 -114 5019 -80
rect 6587 -114 6603 -80
rect 5003 -130 6603 -114
rect 6661 -80 8261 -42
rect 6661 -114 6677 -80
rect 8245 -114 8261 -80
rect 6661 -130 8261 -114
rect 8319 -80 9919 -42
rect 8319 -114 8335 -80
rect 9903 -114 9919 -80
rect 8319 -130 9919 -114
rect 9977 -80 11577 -42
rect 9977 -114 9993 -80
rect 11561 -114 11577 -80
rect 9977 -130 11577 -114
rect 11635 -80 13235 -42
rect 11635 -114 11651 -80
rect 13219 -114 13235 -80
rect 11635 -130 13235 -114
<< polycont >>
rect -13219 80 -11651 114
rect -11561 80 -9993 114
rect -9903 80 -8335 114
rect -8245 80 -6677 114
rect -6587 80 -5019 114
rect -4929 80 -3361 114
rect -3271 80 -1703 114
rect -1613 80 -45 114
rect 45 80 1613 114
rect 1703 80 3271 114
rect 3361 80 4929 114
rect 5019 80 6587 114
rect 6677 80 8245 114
rect 8335 80 9903 114
rect 9993 80 11561 114
rect 11651 80 13219 114
rect -13219 -114 -11651 -80
rect -11561 -114 -9993 -80
rect -9903 -114 -8335 -80
rect -8245 -114 -6677 -80
rect -6587 -114 -5019 -80
rect -4929 -114 -3361 -80
rect -3271 -114 -1703 -80
rect -1613 -114 -45 -80
rect 45 -114 1613 -80
rect 1703 -114 3271 -80
rect 3361 -114 4929 -80
rect 5019 -114 6587 -80
rect 6677 -114 8245 -80
rect 8335 -114 9903 -80
rect 9993 -114 11561 -80
rect 11651 -114 13219 -80
<< locali >>
rect -13415 218 -13319 252
rect 13319 218 13415 252
rect -13415 156 -13381 218
rect 13381 156 13415 218
rect -13235 80 -13219 114
rect -11651 80 -11635 114
rect -11577 80 -11561 114
rect -9993 80 -9977 114
rect -9919 80 -9903 114
rect -8335 80 -8319 114
rect -8261 80 -8245 114
rect -6677 80 -6661 114
rect -6603 80 -6587 114
rect -5019 80 -5003 114
rect -4945 80 -4929 114
rect -3361 80 -3345 114
rect -3287 80 -3271 114
rect -1703 80 -1687 114
rect -1629 80 -1613 114
rect -45 80 -29 114
rect 29 80 45 114
rect 1613 80 1629 114
rect 1687 80 1703 114
rect 3271 80 3287 114
rect 3345 80 3361 114
rect 4929 80 4945 114
rect 5003 80 5019 114
rect 6587 80 6603 114
rect 6661 80 6677 114
rect 8245 80 8261 114
rect 8319 80 8335 114
rect 9903 80 9919 114
rect 9977 80 9993 114
rect 11561 80 11577 114
rect 11635 80 11651 114
rect 13219 80 13235 114
rect -13281 30 -13247 46
rect -13281 -46 -13247 -30
rect -11623 30 -11589 46
rect -11623 -46 -11589 -30
rect -9965 30 -9931 46
rect -9965 -46 -9931 -30
rect -8307 30 -8273 46
rect -8307 -46 -8273 -30
rect -6649 30 -6615 46
rect -6649 -46 -6615 -30
rect -4991 30 -4957 46
rect -4991 -46 -4957 -30
rect -3333 30 -3299 46
rect -3333 -46 -3299 -30
rect -1675 30 -1641 46
rect -1675 -46 -1641 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 1641 30 1675 46
rect 1641 -46 1675 -30
rect 3299 30 3333 46
rect 3299 -46 3333 -30
rect 4957 30 4991 46
rect 4957 -46 4991 -30
rect 6615 30 6649 46
rect 6615 -46 6649 -30
rect 8273 30 8307 46
rect 8273 -46 8307 -30
rect 9931 30 9965 46
rect 9931 -46 9965 -30
rect 11589 30 11623 46
rect 11589 -46 11623 -30
rect 13247 30 13281 46
rect 13247 -46 13281 -30
rect -13235 -114 -13219 -80
rect -11651 -114 -11635 -80
rect -11577 -114 -11561 -80
rect -9993 -114 -9977 -80
rect -9919 -114 -9903 -80
rect -8335 -114 -8319 -80
rect -8261 -114 -8245 -80
rect -6677 -114 -6661 -80
rect -6603 -114 -6587 -80
rect -5019 -114 -5003 -80
rect -4945 -114 -4929 -80
rect -3361 -114 -3345 -80
rect -3287 -114 -3271 -80
rect -1703 -114 -1687 -80
rect -1629 -114 -1613 -80
rect -45 -114 -29 -80
rect 29 -114 45 -80
rect 1613 -114 1629 -80
rect 1687 -114 1703 -80
rect 3271 -114 3287 -80
rect 3345 -114 3361 -80
rect 4929 -114 4945 -80
rect 5003 -114 5019 -80
rect 6587 -114 6603 -80
rect 6661 -114 6677 -80
rect 8245 -114 8261 -80
rect 8319 -114 8335 -80
rect 9903 -114 9919 -80
rect 9977 -114 9993 -80
rect 11561 -114 11577 -80
rect 11635 -114 11651 -80
rect 13219 -114 13235 -80
rect -13415 -218 -13381 -156
rect 13381 -218 13415 -156
rect -13415 -252 -13319 -218
rect 13319 -252 13415 -218
<< viali >>
rect -13219 80 -11651 114
rect -11561 80 -9993 114
rect -9903 80 -8335 114
rect -8245 80 -6677 114
rect -6587 80 -5019 114
rect -4929 80 -3361 114
rect -3271 80 -1703 114
rect -1613 80 -45 114
rect 45 80 1613 114
rect 1703 80 3271 114
rect 3361 80 4929 114
rect 5019 80 6587 114
rect 6677 80 8245 114
rect 8335 80 9903 114
rect 9993 80 11561 114
rect 11651 80 13219 114
rect -13281 -30 -13247 30
rect -11623 -30 -11589 30
rect -9965 -30 -9931 30
rect -8307 -30 -8273 30
rect -6649 -30 -6615 30
rect -4991 -30 -4957 30
rect -3333 -30 -3299 30
rect -1675 -30 -1641 30
rect -17 -30 17 30
rect 1641 -30 1675 30
rect 3299 -30 3333 30
rect 4957 -30 4991 30
rect 6615 -30 6649 30
rect 8273 -30 8307 30
rect 9931 -30 9965 30
rect 11589 -30 11623 30
rect 13247 -30 13281 30
rect -13219 -114 -11651 -80
rect -11561 -114 -9993 -80
rect -9903 -114 -8335 -80
rect -8245 -114 -6677 -80
rect -6587 -114 -5019 -80
rect -4929 -114 -3361 -80
rect -3271 -114 -1703 -80
rect -1613 -114 -45 -80
rect 45 -114 1613 -80
rect 1703 -114 3271 -80
rect 3361 -114 4929 -80
rect 5019 -114 6587 -80
rect 6677 -114 8245 -80
rect 8335 -114 9903 -80
rect 9993 -114 11561 -80
rect 11651 -114 13219 -80
<< metal1 >>
rect -13231 114 -11639 120
rect -13231 80 -13219 114
rect -11651 80 -11639 114
rect -13231 74 -11639 80
rect -11573 114 -9981 120
rect -11573 80 -11561 114
rect -9993 80 -9981 114
rect -11573 74 -9981 80
rect -9915 114 -8323 120
rect -9915 80 -9903 114
rect -8335 80 -8323 114
rect -9915 74 -8323 80
rect -8257 114 -6665 120
rect -8257 80 -8245 114
rect -6677 80 -6665 114
rect -8257 74 -6665 80
rect -6599 114 -5007 120
rect -6599 80 -6587 114
rect -5019 80 -5007 114
rect -6599 74 -5007 80
rect -4941 114 -3349 120
rect -4941 80 -4929 114
rect -3361 80 -3349 114
rect -4941 74 -3349 80
rect -3283 114 -1691 120
rect -3283 80 -3271 114
rect -1703 80 -1691 114
rect -3283 74 -1691 80
rect -1625 114 -33 120
rect -1625 80 -1613 114
rect -45 80 -33 114
rect -1625 74 -33 80
rect 33 114 1625 120
rect 33 80 45 114
rect 1613 80 1625 114
rect 33 74 1625 80
rect 1691 114 3283 120
rect 1691 80 1703 114
rect 3271 80 3283 114
rect 1691 74 3283 80
rect 3349 114 4941 120
rect 3349 80 3361 114
rect 4929 80 4941 114
rect 3349 74 4941 80
rect 5007 114 6599 120
rect 5007 80 5019 114
rect 6587 80 6599 114
rect 5007 74 6599 80
rect 6665 114 8257 120
rect 6665 80 6677 114
rect 8245 80 8257 114
rect 6665 74 8257 80
rect 8323 114 9915 120
rect 8323 80 8335 114
rect 9903 80 9915 114
rect 8323 74 9915 80
rect 9981 114 11573 120
rect 9981 80 9993 114
rect 11561 80 11573 114
rect 9981 74 11573 80
rect 11639 114 13231 120
rect 11639 80 11651 114
rect 13219 80 13231 114
rect 11639 74 13231 80
rect -13287 30 -13241 42
rect -13287 -30 -13281 30
rect -13247 -30 -13241 30
rect -13287 -42 -13241 -30
rect -11629 30 -11583 42
rect -11629 -30 -11623 30
rect -11589 -30 -11583 30
rect -11629 -42 -11583 -30
rect -9971 30 -9925 42
rect -9971 -30 -9965 30
rect -9931 -30 -9925 30
rect -9971 -42 -9925 -30
rect -8313 30 -8267 42
rect -8313 -30 -8307 30
rect -8273 -30 -8267 30
rect -8313 -42 -8267 -30
rect -6655 30 -6609 42
rect -6655 -30 -6649 30
rect -6615 -30 -6609 30
rect -6655 -42 -6609 -30
rect -4997 30 -4951 42
rect -4997 -30 -4991 30
rect -4957 -30 -4951 30
rect -4997 -42 -4951 -30
rect -3339 30 -3293 42
rect -3339 -30 -3333 30
rect -3299 -30 -3293 30
rect -3339 -42 -3293 -30
rect -1681 30 -1635 42
rect -1681 -30 -1675 30
rect -1641 -30 -1635 30
rect -1681 -42 -1635 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 1635 30 1681 42
rect 1635 -30 1641 30
rect 1675 -30 1681 30
rect 1635 -42 1681 -30
rect 3293 30 3339 42
rect 3293 -30 3299 30
rect 3333 -30 3339 30
rect 3293 -42 3339 -30
rect 4951 30 4997 42
rect 4951 -30 4957 30
rect 4991 -30 4997 30
rect 4951 -42 4997 -30
rect 6609 30 6655 42
rect 6609 -30 6615 30
rect 6649 -30 6655 30
rect 6609 -42 6655 -30
rect 8267 30 8313 42
rect 8267 -30 8273 30
rect 8307 -30 8313 30
rect 8267 -42 8313 -30
rect 9925 30 9971 42
rect 9925 -30 9931 30
rect 9965 -30 9971 30
rect 9925 -42 9971 -30
rect 11583 30 11629 42
rect 11583 -30 11589 30
rect 11623 -30 11629 30
rect 11583 -42 11629 -30
rect 13241 30 13287 42
rect 13241 -30 13247 30
rect 13281 -30 13287 30
rect 13241 -42 13287 -30
rect -13231 -80 -11639 -74
rect -13231 -114 -13219 -80
rect -11651 -114 -11639 -80
rect -13231 -120 -11639 -114
rect -11573 -80 -9981 -74
rect -11573 -114 -11561 -80
rect -9993 -114 -9981 -80
rect -11573 -120 -9981 -114
rect -9915 -80 -8323 -74
rect -9915 -114 -9903 -80
rect -8335 -114 -8323 -80
rect -9915 -120 -8323 -114
rect -8257 -80 -6665 -74
rect -8257 -114 -8245 -80
rect -6677 -114 -6665 -80
rect -8257 -120 -6665 -114
rect -6599 -80 -5007 -74
rect -6599 -114 -6587 -80
rect -5019 -114 -5007 -80
rect -6599 -120 -5007 -114
rect -4941 -80 -3349 -74
rect -4941 -114 -4929 -80
rect -3361 -114 -3349 -80
rect -4941 -120 -3349 -114
rect -3283 -80 -1691 -74
rect -3283 -114 -3271 -80
rect -1703 -114 -1691 -80
rect -3283 -120 -1691 -114
rect -1625 -80 -33 -74
rect -1625 -114 -1613 -80
rect -45 -114 -33 -80
rect -1625 -120 -33 -114
rect 33 -80 1625 -74
rect 33 -114 45 -80
rect 1613 -114 1625 -80
rect 33 -120 1625 -114
rect 1691 -80 3283 -74
rect 1691 -114 1703 -80
rect 3271 -114 3283 -80
rect 1691 -120 3283 -114
rect 3349 -80 4941 -74
rect 3349 -114 3361 -80
rect 4929 -114 4941 -80
rect 3349 -120 4941 -114
rect 5007 -80 6599 -74
rect 5007 -114 5019 -80
rect 6587 -114 6599 -80
rect 5007 -120 6599 -114
rect 6665 -80 8257 -74
rect 6665 -114 6677 -80
rect 8245 -114 8257 -80
rect 6665 -120 8257 -114
rect 8323 -80 9915 -74
rect 8323 -114 8335 -80
rect 9903 -114 9915 -80
rect 8323 -120 9915 -114
rect 9981 -80 11573 -74
rect 9981 -114 9993 -80
rect 11561 -114 11573 -80
rect 9981 -120 11573 -114
rect 11639 -80 13231 -74
rect 11639 -114 11651 -80
rect 13219 -114 13231 -80
rect 11639 -120 13231 -114
<< properties >>
string FIXED_BBOX -13398 -235 13398 235
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 8.0 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
