** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/cace/trip_up_down.sch
**.subckt trip_up_down
Vavss avss GND DC 0
Vena ena GND DC 1.8
Vavdd avdd GND pwl (0 2 3m 6 6m 2) DC 3.3
.save i(vavdd)
Vbg1v2 vbg_1v2 GND DC 1.2
Ibias vbp avss 200n
XM1 ibg_200n vbp avdd_bg avdd_bg sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM0 vbp vbp avdd_bg avdd_bg sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vdvss dvss GND DC 0
Vdvdd dvdd GND DC 1.8
.save i(vdvdd)
rsns itest GND 1e6 m=1
cload ovout GND 2e-11 m=1
xIovr avdd avss dvdd dvss vbg_1v2 ovout itest otrip[3] otrip[2] otrip[1] otrip[0] vin ena isrc_sel ibg_200n  sky130_ajc_ip__overvoltage
Vvotrip0 otrip[0] GND DC 0.0
.save i(vvotrip0)
Vvotrip1 otrip[1] GND DC 0.0
.save i(vvotrip1)
Vvotrip2 otrip[2] GND DC 0.0
.save i(vvotrip2)
Vvotrip3 otrip[3] GND DC 1.8
.save i(vvotrip3)
Visrc_sel isrc_sel GND DC 0.0
Vavdd_bg avdd_bg GND DC 3.3
**** begin user architecture code

* CACE gensim simulation file hysteresis_8
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find trip voltage by ramping Vavdd, both up and down.

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
*.include ./netlist/schematic/sky130_ajc_ip__overvoltage.spice


.option TEMP=85
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1
*.option reltol=5e-5
.option reltol=1e-3
.option abstol=1e-3

.save all



.csparam dvdd2=0.9
.control
tran 10u 6m
meas tran vtrip_r find v(avdd) when v(ovout)=$&dvdd2 td=300u rise=1
meas tran vtrip_f find v(avdd) when v(ovout)=$&dvdd2 td=3m fall=1
*meas tran vtrip_r find v(avdd) when v(xiovr.xiana.vl)=$&dvdd2 td=300u rise=1
*meas tran vtrip_f find v(avdd) when v(xiovr.xiana.vl)=$&dvdd2 td=3m fall=1
echo $&vtrip_r > ngspice/hysteresis_8.data
echo $&vtrip_f >> ngspice/hysteresis_8.data
quit
.endc


**** end user architecture code
**.ends

* expanding   symbol:  xschem/sky130_ajc_ip__overvoltage.sym # of pins=12
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/sky130_ajc_ip__overvoltage.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/sky130_ajc_ip__overvoltage.sch
.subckt sky130_ajc_ip__overvoltage avdd avss dvdd dvss vbg_1v2 ovout itest otrip[3] otrip[2] otrip[1] otrip[0] vin ena isrc_sel ibg_200n
*.ipin avdd
*.ipin avss
*.ipin dvdd
*.ipin dvss
*.ipin vbg_1v2
*.ipin otrip[3],otrip[2],otrip[1],otrip[0]
*.ipin ena
*.ipin isrc_sel
*.ipin ibg_200n
*.opin vin
*.opin ovout
*.opin itest
xIana otrip_decoded_15_ otrip_decoded_14_ otrip_decoded_13_ otrip_decoded_12_ otrip_decoded_11_ otrip_decoded_10_ otrip_decoded_9_ otrip_decoded_8_ otrip_decoded_7_ otrip_decoded_6_ otrip_decoded_5_ otrip_decoded_4_ otrip_decoded_3_ otrip_decoded_2_ otrip_decoded_1_ otrip_decoded_0_ vbg_1v2 ena avdd avss dvdd isrc_sel dvss vin itest ibg_200n ovout overvoltage_ana_rcx
**** begin user architecture code



*XSPICE CO-SIM netlist
.include overvoltage_dig.out.spice

r0 otrip[0] otrip0 1
r1 otrip[1] otrip1 1
r2 otrip[2] otrip2 1
r3 otrip[3] otrip3 1

xiovervoltage_dig dvss dvdd otrip0 otrip1 otrip2 otrip3 otrip_decoded_0_ otrip_decoded_10_ otrip_decoded_11_ otrip_decoded_12_ otrip_decoded_13_ otrip_decoded_14_ otrip_decoded_15_ otrip_decoded_1_ otrip_decoded_2_ otrip_decoded_3_ otrip_decoded_4_ otrip_decoded_5_ otrip_decoded_6_ otrip_decoded_7_ otrip_decoded_8_ otrip_decoded_9_ overvoltage_dig



**** end user architecture code
.ends


* expanding   symbol:  xschem/overvoltage_ana_rcx.sym # of pins=12
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/overvoltage_ana_rcx.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/overvoltage_ana_rcx.sch
.subckt overvoltage_ana_rcx otrip_decoded[15] otrip_decoded[14] otrip_decoded[13] otrip_decoded[12] otrip_decoded[11] otrip_decoded[10] otrip_decoded[9] otrip_decoded[8] otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[4] otrip_decoded[3] otrip_decoded[2] otrip_decoded[1] otrip_decoded[0] vbg_1v2 ena avdd avss dvdd isrc_sel dvss vin itest ibg_200n ovout
*.ipin vbg_1v2
*.ipin avdd
*.ipin avss
*.ipin dvdd
*.ipin dvss
*.ipin ena
*.ipin isrc_sel
*.ipin ibg_200n
*.opin ovout
*.opin itest
*.ipin otrip_decoded[15],otrip_decoded[14],otrip_decoded[13],otrip_decoded[12],otrip_decoded[11],otrip_decoded[10],otrip_decoded[9],otrip_decoded[8],otrip_decoded[7],otrip_decoded[6],otrip_decoded[5],otrip_decoded[4],otrip_decoded[3],otrip_decoded[2],otrip_decoded[1],otrip_decoded[0]
*.opin vin
**** begin user architecture code



.include mag/rcx/overvoltage_ana_rcx.spice

xIana otrip_decoded[14] otrip_decoded[13] otrip_decoded[11]  otrip_decoded[10] otrip_decoded[1] otrip_decoded[0] ena itest ibg_200n otrip_decoded[7]  otrip_decoded[4] vbg_1v2 vin isrc_sel otrip_decoded[5] otrip_decoded[8] otrip_decoded[2]  ovout otrip_decoded[15] otrip_decoded[9] otrip_decoded[12] otrip_decoded[3] otrip_decoded[6]  avss dvdd dvss avdd overvoltage_ana_rcx


**** end user architecture code
.ends

.GLOBAL GND
.end
