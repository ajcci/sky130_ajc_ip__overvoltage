magic
tech sky130A
magscale 1 2
timestamp 1712718737
<< error_s >>
rect 26332 18112 26944 22475
rect 27232 22276 27278 22809
rect 26978 21754 27024 22008
rect 27232 21188 27278 21754
rect 26978 20666 27024 20920
rect 27232 20100 27278 20666
rect 26978 19578 27024 19832
rect 27232 19012 27278 19578
<< metal1 >>
rect 573 27559 579 27959
rect 979 27559 985 27959
rect 38495 11718 41643 12028
rect 41953 11718 41959 12028
rect 38553 11462 42086 11662
rect 42286 11462 42292 11662
rect 38481 11206 40724 11406
rect 40924 11206 40930 11406
<< via1 >>
rect 579 27559 979 27959
rect 41643 11718 41953 12028
rect 42086 11462 42286 11662
rect 40724 11206 40924 11406
<< metal2 >>
rect 579 27959 979 27965
rect 123 27494 523 27503
rect 123 25701 523 27094
rect 579 25705 979 27559
rect 8831 21182 8883 28879
rect 9797 21381 9857 28879
rect 10854 16753 10928 28879
rect 13054 13951 13118 28879
rect 25007 27689 25108 27698
rect 25007 26676 25108 27588
rect 37664 23473 37720 23480
rect 26260 23464 26324 23473
rect 22447 20766 22503 20773
rect 22445 20764 22505 20766
rect 22445 20708 22447 20764
rect 22503 20708 22505 20764
rect 20145 18358 20209 18362
rect 20140 18302 20149 18358
rect 20205 18302 20214 18358
rect 13054 13887 13154 13951
rect 13090 13778 13154 13887
rect 20145 13760 20209 18302
rect 20342 15399 20398 15406
rect 20340 15397 20400 15399
rect 20340 15341 20342 15397
rect 20398 15341 20400 15397
rect 20340 13974 20400 15341
rect 22445 13943 22505 20708
rect 24716 16553 24772 16560
rect 24714 16551 24774 16553
rect 24714 16495 24716 16551
rect 24772 16495 24774 16551
rect 24562 15905 24626 15914
rect 22612 15552 22668 15559
rect 22610 15550 22670 15552
rect 22610 15494 22612 15550
rect 22668 15494 22670 15550
rect 22610 13806 22670 15494
rect 24562 13881 24626 15841
rect 20145 13696 20396 13760
rect 20332 12238 20396 13696
rect 22453 13746 22670 13806
rect 24714 13765 24774 16495
rect 25328 16329 25337 16389
rect 25397 16329 25406 16389
rect 26260 15726 26324 23400
rect 37662 23471 37722 23473
rect 37662 23415 37664 23471
rect 37720 23415 37722 23471
rect 37502 22793 37558 22800
rect 37500 22791 37560 22793
rect 26419 22772 26483 22781
rect 26419 15901 26483 22708
rect 37500 22735 37502 22791
rect 37558 22735 37560 22791
rect 37361 22113 37417 22120
rect 37359 22111 37419 22113
rect 26672 22093 26736 22102
rect 26419 15845 26423 15901
rect 26479 15845 26483 15901
rect 26419 15841 26483 15845
rect 26541 21406 26605 21415
rect 26423 15836 26479 15841
rect 26260 15670 26264 15726
rect 26320 15670 26324 15726
rect 26260 15666 26324 15670
rect 26264 15661 26320 15666
rect 22453 12228 22513 13746
rect 24570 13705 24774 13765
rect 26541 13756 26605 21342
rect 26672 18506 26736 22029
rect 37359 22055 37361 22111
rect 37417 22055 37419 22111
rect 36822 21433 36878 21440
rect 36820 21431 36880 21433
rect 36820 21375 36822 21431
rect 36878 21375 36880 21431
rect 26672 18450 26676 18506
rect 26732 18450 26736 18506
rect 26672 18446 26736 18450
rect 32805 18510 32869 18519
rect 26676 18441 26732 18446
rect 30905 18200 30961 18207
rect 30903 18198 30963 18200
rect 30903 18142 30905 18198
rect 30961 18142 30963 18198
rect 28942 17765 28998 17772
rect 28940 17763 29000 17765
rect 28940 17707 28942 17763
rect 28998 17707 29000 17763
rect 26684 17624 26740 17631
rect 26682 17622 26742 17624
rect 26682 17566 26684 17622
rect 26740 17566 26742 17622
rect 26682 14012 26742 17566
rect 28801 15263 28857 15270
rect 28799 15261 28859 15263
rect 28799 15205 28801 15261
rect 28857 15205 28859 15261
rect 28799 13965 28859 15205
rect 28940 13780 29000 17707
rect 30048 15561 30104 16631
rect 30692 16562 30748 16631
rect 30690 16553 30750 16562
rect 30690 16484 30750 16493
rect 30722 15730 30786 15739
rect 30046 15552 30106 15561
rect 30046 15483 30106 15492
rect 24570 12218 24630 13705
rect 26541 13692 26738 13756
rect 26674 12147 26738 13692
rect 28791 13720 29000 13780
rect 30722 13804 30786 15666
rect 30903 13987 30963 18142
rect 31336 15408 31392 16631
rect 31334 15399 31394 15408
rect 31334 15330 31394 15339
rect 31980 15272 32036 16631
rect 32624 15756 32680 16631
rect 32622 15747 32682 15756
rect 32622 15678 32682 15687
rect 31978 15263 32038 15272
rect 31978 15194 32038 15203
rect 30722 13740 30962 13804
rect 28791 12233 28851 13720
rect 30898 12147 30962 13740
rect 32805 13753 32869 18446
rect 35126 18069 35182 18076
rect 35124 18067 35184 18069
rect 35124 18011 35126 18067
rect 35182 18011 35184 18067
rect 33015 17904 33071 17911
rect 33013 17902 33073 17904
rect 33013 17846 33015 17902
rect 33071 17846 33073 17902
rect 33013 13975 33073 17846
rect 33743 16877 33803 16886
rect 33268 16004 33324 16640
rect 33743 16387 33803 16817
rect 33736 16331 33745 16387
rect 33801 16331 33810 16387
rect 33743 16329 33803 16331
rect 33912 16288 33968 16657
rect 34556 16570 34612 16647
rect 34554 16561 34614 16570
rect 34554 16492 34614 16501
rect 33910 16279 33970 16288
rect 33910 16210 33970 16219
rect 33266 15995 33326 16004
rect 33266 15926 33326 15935
rect 35124 13950 35184 18011
rect 36820 17909 36880 21375
rect 36963 20753 37019 20760
rect 36961 20751 37021 20753
rect 36961 20695 36963 20751
rect 37019 20695 37021 20751
rect 36961 18069 37021 20695
rect 37097 20071 37157 20073
rect 37090 20015 37099 20071
rect 37155 20015 37164 20071
rect 37097 19563 37157 20015
rect 37097 19503 37283 19563
rect 37097 19391 37161 19395
rect 37092 19335 37101 19391
rect 37157 19335 37166 19391
rect 37097 18362 37161 19335
rect 37097 18289 37161 18298
rect 37223 18200 37283 19503
rect 37223 18131 37283 18140
rect 36961 18000 37021 18009
rect 36811 17904 36889 17909
rect 36811 17844 36820 17904
rect 36880 17844 36889 17904
rect 36811 17835 36889 17844
rect 37359 17765 37419 22055
rect 37359 17696 37419 17705
rect 37500 17624 37560 22735
rect 37500 17555 37560 17564
rect 35327 17467 35383 17474
rect 37662 17467 37722 23415
rect 35325 17465 35385 17467
rect 35325 17409 35327 17465
rect 35383 17409 35385 17465
rect 35325 13812 35385 17409
rect 37662 17398 37722 17407
rect 37225 13947 37307 13952
rect 37225 13883 37234 13947
rect 37298 13883 37307 13947
rect 37225 13875 37307 13883
rect 32805 13689 33074 13753
rect 33010 12151 33074 13689
rect 35131 13752 35385 13812
rect 35131 12271 35191 13752
rect 37225 12147 37234 12211
rect 37298 12147 37307 12211
rect 41632 12028 41964 12039
rect 41632 11718 41643 12028
rect 41953 11718 41964 12028
rect 41632 11707 41964 11718
rect 42077 11662 42295 11671
rect 42077 11462 42086 11662
rect 42286 11462 42295 11662
rect 42077 11453 42295 11462
rect 40715 11406 40933 11415
rect 40715 11206 40724 11406
rect 40924 11206 40933 11406
rect 40715 11197 40933 11206
rect 582 8086 972 8095
rect 582 7687 972 7696
rect 8809 -1091 9111 5783
rect 9164 -643 9466 5444
rect 9164 -954 9466 -945
rect 8809 -1402 9111 -1393
<< via2 >>
rect 123 27094 523 27494
rect 25007 27588 25108 27689
rect 26260 23400 26324 23464
rect 22447 20708 22503 20764
rect 20149 18302 20205 18358
rect 20342 15341 20398 15397
rect 24716 16495 24772 16551
rect 24562 15841 24626 15905
rect 22612 15494 22668 15550
rect 25337 16329 25397 16389
rect 37664 23415 37720 23471
rect 26419 22708 26483 22772
rect 37502 22735 37558 22791
rect 26672 22029 26736 22093
rect 26423 15845 26479 15901
rect 26541 21342 26605 21406
rect 26264 15670 26320 15726
rect 37361 22055 37417 22111
rect 36822 21375 36878 21431
rect 26676 18450 26732 18506
rect 32805 18446 32869 18510
rect 30905 18142 30961 18198
rect 28942 17707 28998 17763
rect 26684 17566 26740 17622
rect 28801 15205 28857 15261
rect 30690 16493 30750 16553
rect 30722 15666 30786 15730
rect 30046 15492 30106 15552
rect 31334 15339 31394 15399
rect 32622 15687 32682 15747
rect 31978 15203 32038 15263
rect 35126 18011 35182 18067
rect 33015 17846 33071 17902
rect 33743 16817 33803 16877
rect 33745 16331 33801 16387
rect 34554 16501 34614 16561
rect 33910 16219 33970 16279
rect 33266 15935 33326 15995
rect 36963 20695 37019 20751
rect 37099 20015 37155 20071
rect 37101 19335 37157 19391
rect 37097 18298 37161 18362
rect 37223 18140 37283 18200
rect 36961 18009 37021 18069
rect 36820 17844 36880 17904
rect 37359 17705 37419 17765
rect 37500 17564 37560 17624
rect 35327 17409 35383 17465
rect 37662 17407 37722 17467
rect 37234 13883 37298 13947
rect 37234 12147 37298 12211
rect 41643 11718 41953 12028
rect 42086 11462 42286 11662
rect 40724 11206 40924 11406
rect 582 7696 972 8086
rect 123 6835 523 7235
rect 9164 -945 9466 -643
rect 8809 -1393 9111 -1091
<< metal3 >>
rect -2433 28873 42464 28879
rect -2433 28485 -2427 28873
rect -2039 28806 42070 28873
rect -2039 28798 33111 28806
rect -2039 28485 28111 28798
rect -2433 28480 28111 28485
rect 28429 28488 33111 28798
rect 33429 28488 42070 28806
rect 28429 28485 42070 28488
rect 42458 28485 42464 28873
rect 28429 28480 42464 28485
rect -2433 28479 42464 28480
rect -2433 28413 42464 28419
rect -2433 28025 -1967 28413
rect -1579 28373 41610 28413
rect -1579 28055 28771 28373
rect 29089 28356 41610 28373
rect 29089 28055 33771 28356
rect -1579 28038 33771 28055
rect 34089 28038 41610 28356
rect -1579 28025 41610 28038
rect 41998 28025 42464 28413
rect -2433 28019 42464 28025
rect -2433 27953 42464 27959
rect -2433 27565 -1507 27953
rect -1119 27689 41150 27953
rect -1119 27588 25007 27689
rect 25108 27588 41150 27689
rect -1119 27565 41150 27588
rect 41538 27565 42464 27953
rect -2433 27559 42464 27565
rect -2433 27494 42464 27499
rect -2433 27493 123 27494
rect -2433 27105 -1047 27493
rect -659 27105 123 27493
rect -2433 27099 123 27105
rect 118 27094 123 27099
rect 523 27493 42464 27494
rect 523 27105 40690 27493
rect 41078 27105 42464 27493
rect 523 27099 42464 27105
rect 523 27094 528 27099
rect 118 27089 528 27094
rect 37659 23473 37725 23476
rect 37297 23471 37725 23473
rect 26255 23464 26329 23469
rect 26255 23400 26260 23464
rect 26324 23400 26329 23464
rect 37297 23415 37664 23471
rect 37720 23415 37725 23471
rect 37297 23413 37725 23415
rect 37659 23410 37725 23413
rect 26255 23395 26329 23400
rect 37497 22793 37563 22796
rect 37279 22791 37563 22793
rect 26414 22772 26488 22777
rect 26414 22708 26419 22772
rect 26483 22708 26488 22772
rect 37279 22735 37502 22791
rect 37558 22735 37563 22791
rect 37279 22733 37563 22735
rect 37497 22730 37563 22733
rect 26414 22703 26488 22708
rect 37356 22113 37422 22116
rect 37132 22111 37422 22113
rect 26667 22093 26741 22098
rect 26667 22029 26672 22093
rect 26736 22029 26741 22093
rect 37132 22055 37361 22111
rect 37417 22055 37422 22111
rect 37132 22053 37422 22055
rect 37356 22050 37422 22053
rect 26667 22024 26741 22029
rect 36817 21433 36883 21436
rect 36817 21431 37193 21433
rect 26536 21406 26610 21411
rect 26536 21342 26541 21406
rect 26605 21342 26610 21406
rect 36817 21375 36822 21431
rect 36878 21375 37193 21431
rect 36817 21373 37193 21375
rect 36817 21370 36883 21373
rect 26536 21337 26610 21342
rect 22442 20766 22508 20769
rect 22442 20764 26166 20766
rect 22442 20708 22447 20764
rect 22503 20708 26166 20764
rect 22442 20706 26166 20708
rect 36958 20753 37024 20756
rect 36958 20751 37331 20753
rect 22442 20703 22508 20706
rect 36958 20695 36963 20751
rect 37019 20695 37331 20751
rect 36958 20693 37331 20695
rect 36958 20690 37024 20693
rect 37094 20071 37160 20076
rect 37094 20015 37099 20071
rect 37155 20015 37160 20071
rect 37094 20010 37160 20015
rect 37096 19391 37162 19396
rect 37096 19335 37101 19391
rect 37157 19335 37162 19391
rect 37096 19330 37162 19335
rect 26671 18510 26737 18511
rect 32800 18510 32874 18515
rect 26671 18506 32805 18510
rect 26671 18450 26676 18506
rect 26732 18450 32805 18506
rect 26671 18446 32805 18450
rect 32869 18446 32874 18510
rect 26671 18445 26737 18446
rect 32800 18441 32874 18446
rect 20144 18362 20210 18363
rect 37092 18362 37166 18367
rect 20144 18358 37097 18362
rect 20144 18302 20149 18358
rect 20205 18302 37097 18358
rect 20144 18298 37097 18302
rect 37161 18298 37166 18362
rect 20144 18297 20210 18298
rect 37092 18293 37166 18298
rect 30900 18200 30966 18203
rect 37218 18200 37288 18205
rect 30900 18198 37223 18200
rect 30900 18142 30905 18198
rect 30961 18142 37223 18198
rect 30900 18140 37223 18142
rect 37283 18140 37288 18200
rect 30900 18137 30966 18140
rect 37218 18135 37288 18140
rect 35121 18069 35187 18072
rect 36956 18069 37026 18074
rect 35121 18067 36961 18069
rect 35121 18011 35126 18067
rect 35182 18011 36961 18067
rect 35121 18009 36961 18011
rect 37021 18009 37026 18069
rect 35121 18006 35187 18009
rect 36956 18004 37026 18009
rect 33010 17904 33076 17907
rect 36815 17904 36885 17909
rect 33010 17902 36820 17904
rect 33010 17846 33015 17902
rect 33071 17846 36820 17902
rect 33010 17844 36820 17846
rect 36880 17844 36885 17904
rect 33010 17841 33076 17844
rect 36815 17839 36885 17844
rect 28937 17765 29003 17768
rect 37354 17765 37424 17770
rect 28937 17763 37359 17765
rect 28937 17707 28942 17763
rect 28998 17707 37359 17763
rect 28937 17705 37359 17707
rect 37419 17705 37424 17765
rect 28937 17702 29003 17705
rect 37354 17700 37424 17705
rect 26679 17624 26745 17627
rect 37495 17624 37565 17629
rect 26679 17622 37500 17624
rect 26679 17566 26684 17622
rect 26740 17566 37500 17622
rect 26679 17564 37500 17566
rect 37560 17564 37565 17624
rect 26679 17561 26745 17564
rect 37495 17559 37565 17564
rect 35322 17467 35388 17470
rect 37657 17467 37727 17472
rect 35322 17465 37662 17467
rect 35322 17409 35327 17465
rect 35383 17409 37662 17465
rect 35322 17407 37662 17409
rect 37722 17407 37727 17467
rect 35322 17404 35388 17407
rect 37657 17402 37727 17407
rect 33738 16877 33808 16882
rect 33738 16817 33743 16877
rect 33803 16817 42464 16877
rect 33738 16812 33808 16817
rect 34549 16561 34619 16566
rect 24711 16553 24777 16556
rect 30685 16553 30755 16558
rect 24711 16551 30690 16553
rect 24711 16495 24716 16551
rect 24772 16495 30690 16551
rect 24711 16493 30690 16495
rect 30750 16493 30755 16553
rect 34549 16501 34554 16561
rect 34614 16501 42464 16561
rect 34549 16496 34619 16501
rect 24711 16490 24777 16493
rect 30685 16488 30755 16493
rect 25332 16389 25402 16394
rect 33740 16389 33806 16392
rect 25332 16329 25337 16389
rect 25397 16387 33806 16389
rect 25397 16331 33745 16387
rect 33801 16331 33806 16387
rect 25397 16329 33806 16331
rect 25332 16324 25402 16329
rect 33740 16326 33806 16329
rect 33905 16279 33975 16284
rect 33905 16219 33910 16279
rect 33970 16219 42464 16279
rect 33905 16214 33975 16219
rect 33261 15995 33331 16000
rect 33261 15935 33266 15995
rect 33326 15935 42464 15995
rect 33261 15930 33331 15935
rect 24557 15905 24631 15910
rect 26418 15905 26484 15906
rect 24557 15841 24562 15905
rect 24626 15901 26484 15905
rect 24626 15845 26423 15901
rect 26479 15845 26484 15901
rect 24626 15841 26484 15845
rect 24557 15836 24631 15841
rect 26418 15840 26484 15841
rect 32617 15747 32687 15752
rect 26259 15730 26325 15731
rect 30717 15730 30791 15735
rect 26259 15726 30722 15730
rect 26259 15670 26264 15726
rect 26320 15670 30722 15726
rect 26259 15666 30722 15670
rect 30786 15666 30791 15730
rect 32617 15687 32622 15747
rect 32682 15687 42464 15747
rect 32617 15682 32687 15687
rect 26259 15665 26325 15666
rect 30717 15661 30791 15666
rect 22607 15552 22673 15555
rect 30041 15552 30111 15557
rect 22607 15550 30046 15552
rect 22607 15494 22612 15550
rect 22668 15494 30046 15550
rect 22607 15492 30046 15494
rect 30106 15492 30111 15552
rect 22607 15489 22673 15492
rect 30041 15487 30111 15492
rect 20337 15399 20403 15402
rect 31329 15399 31399 15404
rect 20337 15397 31334 15399
rect 20337 15341 20342 15397
rect 20398 15341 31334 15397
rect 20337 15339 31334 15341
rect 31394 15339 31399 15399
rect 20337 15336 20403 15339
rect 31329 15334 31399 15339
rect 28796 15263 28862 15266
rect 31973 15263 32043 15268
rect 28796 15261 31978 15263
rect 28796 15205 28801 15261
rect 28857 15205 31978 15261
rect 28796 15203 31978 15205
rect 32038 15203 32043 15263
rect 28796 15200 28862 15203
rect 31973 15198 32043 15203
rect 4513 14168 4583 14238
rect 37229 13947 37303 13952
rect 37229 13883 37234 13947
rect 37298 13883 42464 13947
rect 37229 13878 37303 13883
rect 37229 12211 37303 12216
rect 37229 12147 37234 12211
rect 37298 12147 42464 12211
rect 37229 12142 37303 12147
rect 41632 12033 41964 12039
rect 41632 11713 41638 12033
rect 41958 11713 41964 12033
rect 41632 11707 41964 11713
rect 42077 11662 42295 11671
rect 42077 11462 42086 11662
rect 42286 11462 42295 11662
rect 42077 11453 42295 11462
rect 40715 11406 40933 11415
rect 40715 11206 40724 11406
rect 40924 11206 40933 11406
rect 40715 11197 40933 11206
rect -1518 8091 -1113 8096
rect -1518 8090 977 8091
rect -1518 7692 -1512 8090
rect -1114 8086 977 8090
rect -1114 7696 582 8086
rect 972 7696 977 8086
rect -1114 7692 977 7696
rect -1518 7691 977 7692
rect -1518 7686 -1113 7691
rect 118 7235 528 7240
rect -1056 6835 -1050 7235
rect -650 6835 123 7235
rect 523 6835 528 7235
rect 118 6830 528 6835
rect -2433 -616 42464 -610
rect -2433 -1004 -1047 -616
rect -659 -643 40690 -616
rect -659 -945 9164 -643
rect 9466 -945 40690 -643
rect -659 -1004 40690 -945
rect 41078 -1004 42464 -616
rect -2433 -1010 42464 -1004
rect -2433 -1076 42464 -1070
rect -2433 -1464 -1507 -1076
rect -1119 -1091 41150 -1076
rect -1119 -1393 8809 -1091
rect 9111 -1393 41150 -1091
rect -1119 -1464 41150 -1393
rect 41538 -1464 42464 -1076
rect -2433 -1470 42464 -1464
rect -2433 -1536 42464 -1530
rect -2433 -1924 -1967 -1536
rect -1579 -1924 41610 -1536
rect 41998 -1924 42464 -1536
rect -2433 -1930 42464 -1924
rect -2433 -1996 42464 -1990
rect -2433 -2384 -2427 -1996
rect -2039 -2384 42070 -1996
rect 42458 -2384 42464 -1996
rect -2433 -2390 42464 -2384
<< via3 >>
rect -2427 28485 -2039 28873
rect 28111 28480 28429 28798
rect 33111 28488 33429 28806
rect 42070 28485 42458 28873
rect -1967 28025 -1579 28413
rect 28771 28055 29089 28373
rect 33771 28038 34089 28356
rect 41610 28025 41998 28413
rect -1507 27565 -1119 27953
rect 41150 27565 41538 27953
rect -1047 27105 -659 27493
rect 40690 27105 41078 27493
rect 41638 12028 41958 12033
rect 41638 11718 41643 12028
rect 41643 11718 41953 12028
rect 41953 11718 41958 12028
rect 41638 11713 41958 11718
rect 42086 11462 42286 11662
rect 40724 11206 40924 11406
rect -1512 7692 -1114 8090
rect -1050 6835 -650 7235
rect -1047 -1004 -659 -616
rect 40690 -1004 41078 -616
rect -1507 -1464 -1119 -1076
rect 41150 -1464 41538 -1076
rect -1967 -1924 -1579 -1536
rect 41610 -1924 41998 -1536
rect -2427 -2384 -2039 -1996
rect 42070 -2384 42458 -1996
<< metal4 >>
rect -2433 28873 -2033 28880
rect -2433 28485 -2427 28873
rect -2039 28485 -2033 28873
rect -2433 -1996 -2033 28485
rect -2433 -2384 -2427 -1996
rect -2039 -2384 -2033 -1996
rect -2433 -2390 -2033 -2384
rect -1973 28413 -1573 28880
rect -1973 28025 -1967 28413
rect -1579 28025 -1573 28413
rect -1973 -1536 -1573 28025
rect -1973 -1924 -1967 -1536
rect -1579 -1924 -1573 -1536
rect -1973 -2390 -1573 -1924
rect -1513 27953 -1113 28880
rect -1513 27565 -1507 27953
rect -1119 27565 -1113 27953
rect -1513 8090 -1113 27565
rect -1513 7692 -1512 8090
rect -1114 7692 -1113 8090
rect -1513 -1076 -1113 7692
rect -1513 -1464 -1507 -1076
rect -1119 -1464 -1113 -1076
rect -1513 -2390 -1113 -1464
rect -1053 27493 -653 28880
rect 33110 28806 33430 28807
rect -1053 27105 -1047 27493
rect -659 27105 -653 27493
rect -1053 7236 -653 27105
rect 28110 28798 28430 28799
rect 28110 28480 28111 28798
rect 28429 28480 28430 28798
rect 28110 26029 28430 28480
rect 33110 28488 33111 28806
rect 33429 28488 33430 28806
rect 28770 28373 29090 28374
rect 28770 28055 28771 28373
rect 29089 28055 29090 28373
rect 28770 25980 29090 28055
rect 33110 26095 33430 28488
rect 33770 28356 34090 28357
rect 33770 28038 33771 28356
rect 34089 28038 34090 28356
rect 33770 26015 34090 28038
rect 40684 27493 41084 28880
rect 40684 27105 40690 27493
rect 41078 27105 41084 27493
rect 40684 11406 41084 27105
rect 40684 11206 40724 11406
rect 40924 11206 41084 11406
rect -1053 7235 -649 7236
rect -1053 6835 -1050 7235
rect -650 6835 -649 7235
rect -1053 6834 -649 6835
rect -1053 -616 -653 6834
rect -1053 -1004 -1047 -616
rect -659 -1004 -653 -616
rect -1053 -2390 -653 -1004
rect 40684 -616 41084 11206
rect 40684 -1004 40690 -616
rect 41078 -1004 41084 -616
rect 40684 -2390 41084 -1004
rect 41144 27953 41544 28880
rect 41144 27565 41150 27953
rect 41538 27565 41544 27953
rect 41144 -1076 41544 27565
rect 41144 -1464 41150 -1076
rect 41538 -1464 41544 -1076
rect 41144 -2390 41544 -1464
rect 41604 28413 42004 28880
rect 41604 28025 41610 28413
rect 41998 28025 42004 28413
rect 41604 20547 42004 28025
rect 41604 20275 41689 20547
rect 41961 20275 42004 20547
rect 41604 12033 42004 20275
rect 41604 11713 41638 12033
rect 41958 11713 42004 12033
rect 41604 -1536 42004 11713
rect 41604 -1924 41610 -1536
rect 41998 -1924 42004 -1536
rect 41604 -2390 42004 -1924
rect 42064 28873 42464 28880
rect 42064 28485 42070 28873
rect 42458 28485 42464 28873
rect 42064 19887 42464 28485
rect 42064 19615 42146 19887
rect 42418 19615 42464 19887
rect 42064 11662 42464 19615
rect 42064 11462 42086 11662
rect 42286 11462 42464 11662
rect 42064 -1996 42464 11462
rect 42064 -2384 42070 -1996
rect 42458 -2384 42464 -1996
rect 42064 -2390 42464 -2384
<< via4 >>
rect 41689 20275 41961 20547
rect 42146 19615 42418 19887
<< metal5 >>
rect 36585 20547 41985 20571
rect 36585 20275 41689 20547
rect 41961 20275 41985 20547
rect 36585 20251 41985 20275
rect 36568 19887 42442 19911
rect 36568 19615 42146 19887
rect 42418 19615 42442 19887
rect 36568 19591 42442 19615
use overvoltage_ana  overvoltage_ana_0
timestamp 1712718737
transform 1 0 28385 0 1 16000
box -29038 -16610 12299 11100
use overvoltage_dig  overvoltage_dig_0
timestamp 1712531369
transform 1 0 26166 0 1 16575
box 0 0 12000 9840
<< labels >>
flabel metal3 894 -1930 894 -1930 0 FreeSans 1600 0 0 0 dvss
port 4 nsew
flabel metal3 894 -1470 894 -1470 0 FreeSans 1600 0 0 0 avss
port 2 nsew
flabel metal3 894 -1010 894 -1010 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal3 42464 15715 42464 15715 0 FreeSans 1280 0 0 0 otrip[0]
port 11 nsew
flabel metal3 42464 15964 42464 15964 0 FreeSans 1280 0 0 0 otrip[1]
port 10 nsew
flabel metal3 42464 16248 42464 16248 0 FreeSans 1280 0 0 0 otrip[2]
port 9 nsew
flabel metal3 42464 16529 42464 16529 0 FreeSans 1280 0 0 0 otrip[3]
port 8 nsew
flabel metal3 42464 16846 42464 16846 0 FreeSans 1280 0 0 0 ovout
port 6 nsew
flabel metal2 10891 28879 10891 28879 0 FreeSans 1280 0 0 0 itest
port 7 nsew
flabel metal2 8857 28879 8857 28879 0 FreeSans 1280 0 0 0 vbg_1v2
port 5 nsew
flabel metal2 9828 28879 9828 28879 0 FreeSans 1280 0 0 0 vin
port 12 nsew
flabel metal3 42464 12177 42464 12177 0 FreeSans 1280 0 0 0 ena
port 13 nsew
flabel metal3 42464 13915 42464 13915 0 FreeSans 1280 0 0 0 isrc_sel
port 14 nsew
flabel metal2 13085 28879 13085 28879 0 FreeSans 1280 0 0 0 ibg_200n
port 15 nsew
flabel metal3 894 -2390 894 -2390 0 FreeSans 1600 0 0 0 dvdd
port 3 nsew
<< end >>
