magic
tech sky130A
magscale 1 2
timestamp 1711774300
<< nwell >>
rect -5203 -362 5203 362
<< mvpmos >>
rect -4945 -64 -3345 136
rect -3287 -64 -1687 136
rect -1629 -64 -29 136
rect 29 -64 1629 136
rect 1687 -64 3287 136
rect 3345 -64 4945 136
<< mvpdiff >>
rect -5003 124 -4945 136
rect -5003 -52 -4991 124
rect -4957 -52 -4945 124
rect -5003 -64 -4945 -52
rect -3345 124 -3287 136
rect -3345 -52 -3333 124
rect -3299 -52 -3287 124
rect -3345 -64 -3287 -52
rect -1687 124 -1629 136
rect -1687 -52 -1675 124
rect -1641 -52 -1629 124
rect -1687 -64 -1629 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 1629 124 1687 136
rect 1629 -52 1641 124
rect 1675 -52 1687 124
rect 1629 -64 1687 -52
rect 3287 124 3345 136
rect 3287 -52 3299 124
rect 3333 -52 3345 124
rect 3287 -64 3345 -52
rect 4945 124 5003 136
rect 4945 -52 4957 124
rect 4991 -52 5003 124
rect 4945 -64 5003 -52
<< mvpdiffc >>
rect -4991 -52 -4957 124
rect -3333 -52 -3299 124
rect -1675 -52 -1641 124
rect -17 -52 17 124
rect 1641 -52 1675 124
rect 3299 -52 3333 124
rect 4957 -52 4991 124
<< mvnsubdiff >>
rect -5137 284 5137 296
rect -5137 250 -5029 284
rect 5029 250 5137 284
rect -5137 238 5137 250
rect -5137 188 -5079 238
rect -5137 -188 -5125 188
rect -5091 -188 -5079 188
rect 5079 188 5137 238
rect -5137 -238 -5079 -188
rect 5079 -188 5091 188
rect 5125 -188 5137 188
rect 5079 -238 5137 -188
rect -5137 -250 5137 -238
rect -5137 -284 -5029 -250
rect 5029 -284 5137 -250
rect -5137 -296 5137 -284
<< mvnsubdiffcont >>
rect -5029 250 5029 284
rect -5125 -188 -5091 188
rect 5091 -188 5125 188
rect -5029 -284 5029 -250
<< poly >>
rect -4945 136 -3345 162
rect -3287 136 -1687 162
rect -1629 136 -29 162
rect 29 136 1629 162
rect 1687 136 3287 162
rect 3345 136 4945 162
rect -4945 -111 -3345 -64
rect -4945 -145 -4929 -111
rect -3361 -145 -3345 -111
rect -4945 -161 -3345 -145
rect -3287 -111 -1687 -64
rect -3287 -145 -3271 -111
rect -1703 -145 -1687 -111
rect -3287 -161 -1687 -145
rect -1629 -111 -29 -64
rect -1629 -145 -1613 -111
rect -45 -145 -29 -111
rect -1629 -161 -29 -145
rect 29 -111 1629 -64
rect 29 -145 45 -111
rect 1613 -145 1629 -111
rect 29 -161 1629 -145
rect 1687 -111 3287 -64
rect 1687 -145 1703 -111
rect 3271 -145 3287 -111
rect 1687 -161 3287 -145
rect 3345 -111 4945 -64
rect 3345 -145 3361 -111
rect 4929 -145 4945 -111
rect 3345 -161 4945 -145
<< polycont >>
rect -4929 -145 -3361 -111
rect -3271 -145 -1703 -111
rect -1613 -145 -45 -111
rect 45 -145 1613 -111
rect 1703 -145 3271 -111
rect 3361 -145 4929 -111
<< locali >>
rect -5125 250 -5029 284
rect 5029 250 5125 284
rect -5125 188 -5091 250
rect 5091 188 5125 250
rect -4991 124 -4957 140
rect -4991 -68 -4957 -52
rect -3333 124 -3299 140
rect -3333 -68 -3299 -52
rect -1675 124 -1641 140
rect -1675 -68 -1641 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 1641 124 1675 140
rect 1641 -68 1675 -52
rect 3299 124 3333 140
rect 3299 -68 3333 -52
rect 4957 124 4991 140
rect 4957 -68 4991 -52
rect -4945 -145 -4929 -111
rect -3361 -145 -3345 -111
rect -3287 -145 -3271 -111
rect -1703 -145 -1687 -111
rect -1629 -145 -1613 -111
rect -45 -145 -29 -111
rect 29 -145 45 -111
rect 1613 -145 1629 -111
rect 1687 -145 1703 -111
rect 3271 -145 3287 -111
rect 3345 -145 3361 -111
rect 4929 -145 4945 -111
rect -5125 -250 -5091 -188
rect 5091 -250 5125 -188
rect -5125 -284 -5029 -250
rect 5029 -284 5125 -250
<< viali >>
rect -4991 -52 -4957 124
rect -3333 -52 -3299 124
rect -1675 -52 -1641 124
rect -17 -52 17 124
rect 1641 -52 1675 124
rect 3299 -52 3333 124
rect 4957 -52 4991 124
rect -4929 -145 -3361 -111
rect -3271 -145 -1703 -111
rect -1613 -145 -45 -111
rect 45 -145 1613 -111
rect 1703 -145 3271 -111
rect 3361 -145 4929 -111
<< metal1 >>
rect -4997 124 -4951 136
rect -4997 -52 -4991 124
rect -4957 -52 -4951 124
rect -4997 -64 -4951 -52
rect -3339 124 -3293 136
rect -3339 -52 -3333 124
rect -3299 -52 -3293 124
rect -3339 -64 -3293 -52
rect -1681 124 -1635 136
rect -1681 -52 -1675 124
rect -1641 -52 -1635 124
rect -1681 -64 -1635 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 1635 124 1681 136
rect 1635 -52 1641 124
rect 1675 -52 1681 124
rect 1635 -64 1681 -52
rect 3293 124 3339 136
rect 3293 -52 3299 124
rect 3333 -52 3339 124
rect 3293 -64 3339 -52
rect 4951 124 4997 136
rect 4951 -52 4957 124
rect 4991 -52 4997 124
rect 4951 -64 4997 -52
rect -4941 -111 -3349 -105
rect -4941 -145 -4929 -111
rect -3361 -145 -3349 -111
rect -4941 -151 -3349 -145
rect -3283 -111 -1691 -105
rect -3283 -145 -3271 -111
rect -1703 -145 -1691 -111
rect -3283 -151 -1691 -145
rect -1625 -111 -33 -105
rect -1625 -145 -1613 -111
rect -45 -145 -33 -111
rect -1625 -151 -33 -145
rect 33 -111 1625 -105
rect 33 -145 45 -111
rect 1613 -145 1625 -111
rect 33 -151 1625 -145
rect 1691 -111 3283 -105
rect 1691 -145 1703 -111
rect 3271 -145 3283 -111
rect 1691 -151 3283 -145
rect 3349 -111 4941 -105
rect 3349 -145 3361 -111
rect 4929 -145 4941 -111
rect 3349 -151 4941 -145
<< properties >>
string FIXED_BBOX -5108 -267 5108 267
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 8 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
