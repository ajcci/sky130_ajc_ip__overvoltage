magic
tech sky130A
magscale 1 2
timestamp 1711636687
<< nwell >>
rect -941 -339 941 339
<< mvpmos >>
rect -683 -42 -563 42
rect -505 -42 -385 42
rect -327 -42 -207 42
rect -149 -42 -29 42
rect 29 -42 149 42
rect 207 -42 327 42
rect 385 -42 505 42
rect 563 -42 683 42
<< mvpdiff >>
rect -741 30 -683 42
rect -741 -30 -729 30
rect -695 -30 -683 30
rect -741 -42 -683 -30
rect -563 30 -505 42
rect -563 -30 -551 30
rect -517 -30 -505 30
rect -563 -42 -505 -30
rect -385 30 -327 42
rect -385 -30 -373 30
rect -339 -30 -327 30
rect -385 -42 -327 -30
rect -207 30 -149 42
rect -207 -30 -195 30
rect -161 -30 -149 30
rect -207 -42 -149 -30
rect -29 30 29 42
rect -29 -30 -17 30
rect 17 -30 29 30
rect -29 -42 29 -30
rect 149 30 207 42
rect 149 -30 161 30
rect 195 -30 207 30
rect 149 -42 207 -30
rect 327 30 385 42
rect 327 -30 339 30
rect 373 -30 385 30
rect 327 -42 385 -30
rect 505 30 563 42
rect 505 -30 517 30
rect 551 -30 563 30
rect 505 -42 563 -30
rect 683 30 741 42
rect 683 -30 695 30
rect 729 -30 741 30
rect 683 -42 741 -30
<< mvpdiffc >>
rect -729 -30 -695 30
rect -551 -30 -517 30
rect -373 -30 -339 30
rect -195 -30 -161 30
rect -17 -30 17 30
rect 161 -30 195 30
rect 339 -30 373 30
rect 517 -30 551 30
rect 695 -30 729 30
<< mvnsubdiff >>
rect -875 261 875 273
rect -875 227 -767 261
rect 767 227 875 261
rect -875 215 875 227
rect -875 165 -817 215
rect -875 -165 -863 165
rect -829 -165 -817 165
rect 817 165 875 215
rect -875 -215 -817 -165
rect 817 -165 829 165
rect 863 -165 875 165
rect 817 -215 875 -165
rect -875 -227 875 -215
rect -875 -261 -767 -227
rect 767 -261 875 -227
rect -875 -273 875 -261
<< mvnsubdiffcont >>
rect -767 227 767 261
rect -863 -165 -829 165
rect 829 -165 863 165
rect -767 -261 767 -227
<< poly >>
rect -683 123 -563 139
rect -683 89 -667 123
rect -579 89 -563 123
rect -683 42 -563 89
rect -505 123 -385 139
rect -505 89 -489 123
rect -401 89 -385 123
rect -505 42 -385 89
rect -327 123 -207 139
rect -327 89 -311 123
rect -223 89 -207 123
rect -327 42 -207 89
rect -149 123 -29 139
rect -149 89 -133 123
rect -45 89 -29 123
rect -149 42 -29 89
rect 29 123 149 139
rect 29 89 45 123
rect 133 89 149 123
rect 29 42 149 89
rect 207 123 327 139
rect 207 89 223 123
rect 311 89 327 123
rect 207 42 327 89
rect 385 123 505 139
rect 385 89 401 123
rect 489 89 505 123
rect 385 42 505 89
rect 563 123 683 139
rect 563 89 579 123
rect 667 89 683 123
rect 563 42 683 89
rect -683 -89 -563 -42
rect -683 -123 -667 -89
rect -579 -123 -563 -89
rect -683 -139 -563 -123
rect -505 -89 -385 -42
rect -505 -123 -489 -89
rect -401 -123 -385 -89
rect -505 -139 -385 -123
rect -327 -89 -207 -42
rect -327 -123 -311 -89
rect -223 -123 -207 -89
rect -327 -139 -207 -123
rect -149 -89 -29 -42
rect -149 -123 -133 -89
rect -45 -123 -29 -89
rect -149 -139 -29 -123
rect 29 -89 149 -42
rect 29 -123 45 -89
rect 133 -123 149 -89
rect 29 -139 149 -123
rect 207 -89 327 -42
rect 207 -123 223 -89
rect 311 -123 327 -89
rect 207 -139 327 -123
rect 385 -89 505 -42
rect 385 -123 401 -89
rect 489 -123 505 -89
rect 385 -139 505 -123
rect 563 -89 683 -42
rect 563 -123 579 -89
rect 667 -123 683 -89
rect 563 -139 683 -123
<< polycont >>
rect -667 89 -579 123
rect -489 89 -401 123
rect -311 89 -223 123
rect -133 89 -45 123
rect 45 89 133 123
rect 223 89 311 123
rect 401 89 489 123
rect 579 89 667 123
rect -667 -123 -579 -89
rect -489 -123 -401 -89
rect -311 -123 -223 -89
rect -133 -123 -45 -89
rect 45 -123 133 -89
rect 223 -123 311 -89
rect 401 -123 489 -89
rect 579 -123 667 -89
<< locali >>
rect -863 227 -767 261
rect 767 227 863 261
rect -863 165 -829 227
rect 829 165 863 227
rect -683 89 -667 123
rect -579 89 -563 123
rect -505 89 -489 123
rect -401 89 -385 123
rect -327 89 -311 123
rect -223 89 -207 123
rect -149 89 -133 123
rect -45 89 -29 123
rect 29 89 45 123
rect 133 89 149 123
rect 207 89 223 123
rect 311 89 327 123
rect 385 89 401 123
rect 489 89 505 123
rect 563 89 579 123
rect 667 89 683 123
rect -729 30 -695 46
rect -729 -46 -695 -30
rect -551 30 -517 46
rect -551 -46 -517 -30
rect -373 30 -339 46
rect -373 -46 -339 -30
rect -195 30 -161 46
rect -195 -46 -161 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 161 30 195 46
rect 161 -46 195 -30
rect 339 30 373 46
rect 339 -46 373 -30
rect 517 30 551 46
rect 517 -46 551 -30
rect 695 30 729 46
rect 695 -46 729 -30
rect -683 -123 -667 -89
rect -579 -123 -563 -89
rect -505 -123 -489 -89
rect -401 -123 -385 -89
rect -327 -123 -311 -89
rect -223 -123 -207 -89
rect -149 -123 -133 -89
rect -45 -123 -29 -89
rect 29 -123 45 -89
rect 133 -123 149 -89
rect 207 -123 223 -89
rect 311 -123 327 -89
rect 385 -123 401 -89
rect 489 -123 505 -89
rect 563 -123 579 -89
rect 667 -123 683 -89
rect -863 -227 -829 -165
rect 829 -227 863 -165
rect -863 -261 -767 -227
rect 767 -261 863 -227
<< viali >>
rect -667 89 -579 123
rect -489 89 -401 123
rect -311 89 -223 123
rect -133 89 -45 123
rect 45 89 133 123
rect 223 89 311 123
rect 401 89 489 123
rect 579 89 667 123
rect -729 -30 -695 30
rect -551 -30 -517 30
rect -373 -30 -339 30
rect -195 -30 -161 30
rect -17 -30 17 30
rect 161 -30 195 30
rect 339 -30 373 30
rect 517 -30 551 30
rect 695 -30 729 30
rect -667 -123 -579 -89
rect -489 -123 -401 -89
rect -311 -123 -223 -89
rect -133 -123 -45 -89
rect 45 -123 133 -89
rect 223 -123 311 -89
rect 401 -123 489 -89
rect 579 -123 667 -89
<< metal1 >>
rect -679 123 -567 129
rect -679 89 -667 123
rect -579 89 -567 123
rect -679 83 -567 89
rect -501 123 -389 129
rect -501 89 -489 123
rect -401 89 -389 123
rect -501 83 -389 89
rect -323 123 -211 129
rect -323 89 -311 123
rect -223 89 -211 123
rect -323 83 -211 89
rect -145 123 -33 129
rect -145 89 -133 123
rect -45 89 -33 123
rect -145 83 -33 89
rect 33 123 145 129
rect 33 89 45 123
rect 133 89 145 123
rect 33 83 145 89
rect 211 123 323 129
rect 211 89 223 123
rect 311 89 323 123
rect 211 83 323 89
rect 389 123 501 129
rect 389 89 401 123
rect 489 89 501 123
rect 389 83 501 89
rect 567 123 679 129
rect 567 89 579 123
rect 667 89 679 123
rect 567 83 679 89
rect -735 30 -689 42
rect -735 -30 -729 30
rect -695 -30 -689 30
rect -735 -42 -689 -30
rect -557 30 -511 42
rect -557 -30 -551 30
rect -517 -30 -511 30
rect -557 -42 -511 -30
rect -379 30 -333 42
rect -379 -30 -373 30
rect -339 -30 -333 30
rect -379 -42 -333 -30
rect -201 30 -155 42
rect -201 -30 -195 30
rect -161 -30 -155 30
rect -201 -42 -155 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 155 30 201 42
rect 155 -30 161 30
rect 195 -30 201 30
rect 155 -42 201 -30
rect 333 30 379 42
rect 333 -30 339 30
rect 373 -30 379 30
rect 333 -42 379 -30
rect 511 30 557 42
rect 511 -30 517 30
rect 551 -30 557 30
rect 511 -42 557 -30
rect 689 30 735 42
rect 689 -30 695 30
rect 729 -30 735 30
rect 689 -42 735 -30
rect -679 -89 -567 -83
rect -679 -123 -667 -89
rect -579 -123 -567 -89
rect -679 -129 -567 -123
rect -501 -89 -389 -83
rect -501 -123 -489 -89
rect -401 -123 -389 -89
rect -501 -129 -389 -123
rect -323 -89 -211 -83
rect -323 -123 -311 -89
rect -223 -123 -211 -89
rect -323 -129 -211 -123
rect -145 -89 -33 -83
rect -145 -123 -133 -89
rect -45 -123 -33 -89
rect -145 -129 -33 -123
rect 33 -89 145 -83
rect 33 -123 45 -89
rect 133 -123 145 -89
rect 33 -129 145 -123
rect 211 -89 323 -83
rect 211 -123 223 -89
rect 311 -123 323 -89
rect 211 -129 323 -123
rect 389 -89 501 -83
rect 389 -123 401 -89
rect 489 -123 501 -89
rect 389 -129 501 -123
rect 567 -89 679 -83
rect 567 -123 579 -89
rect 667 -123 679 -89
rect 567 -129 679 -123
<< properties >>
string FIXED_BBOX -846 -244 846 244
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.6 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
