magic
tech sky130A
magscale 1 2
timestamp 1711596774
<< mvnmos >>
rect -4945 -500 -3345 500
rect -3287 -500 -1687 500
rect -1629 -500 -29 500
rect 29 -500 1629 500
rect 1687 -500 3287 500
rect 3345 -500 4945 500
<< mvndiff >>
rect -5003 488 -4945 500
rect -5003 -488 -4991 488
rect -4957 -488 -4945 488
rect -5003 -500 -4945 -488
rect -3345 488 -3287 500
rect -3345 -488 -3333 488
rect -3299 -488 -3287 488
rect -3345 -500 -3287 -488
rect -1687 488 -1629 500
rect -1687 -488 -1675 488
rect -1641 -488 -1629 488
rect -1687 -500 -1629 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 1629 488 1687 500
rect 1629 -488 1641 488
rect 1675 -488 1687 488
rect 1629 -500 1687 -488
rect 3287 488 3345 500
rect 3287 -488 3299 488
rect 3333 -488 3345 488
rect 3287 -500 3345 -488
rect 4945 488 5003 500
rect 4945 -488 4957 488
rect 4991 -488 5003 488
rect 4945 -500 5003 -488
<< mvndiffc >>
rect -4991 -488 -4957 488
rect -3333 -488 -3299 488
rect -1675 -488 -1641 488
rect -17 -488 17 488
rect 1641 -488 1675 488
rect 3299 -488 3333 488
rect 4957 -488 4991 488
<< poly >>
rect -4945 572 -3345 588
rect -4945 538 -4929 572
rect -3361 538 -3345 572
rect -4945 500 -3345 538
rect -3287 572 -1687 588
rect -3287 538 -3271 572
rect -1703 538 -1687 572
rect -3287 500 -1687 538
rect -1629 572 -29 588
rect -1629 538 -1613 572
rect -45 538 -29 572
rect -1629 500 -29 538
rect 29 572 1629 588
rect 29 538 45 572
rect 1613 538 1629 572
rect 29 500 1629 538
rect 1687 572 3287 588
rect 1687 538 1703 572
rect 3271 538 3287 572
rect 1687 500 3287 538
rect 3345 572 4945 588
rect 3345 538 3361 572
rect 4929 538 4945 572
rect 3345 500 4945 538
rect -4945 -538 -3345 -500
rect -4945 -572 -4929 -538
rect -3361 -572 -3345 -538
rect -4945 -588 -3345 -572
rect -3287 -538 -1687 -500
rect -3287 -572 -3271 -538
rect -1703 -572 -1687 -538
rect -3287 -588 -1687 -572
rect -1629 -538 -29 -500
rect -1629 -572 -1613 -538
rect -45 -572 -29 -538
rect -1629 -588 -29 -572
rect 29 -538 1629 -500
rect 29 -572 45 -538
rect 1613 -572 1629 -538
rect 29 -588 1629 -572
rect 1687 -538 3287 -500
rect 1687 -572 1703 -538
rect 3271 -572 3287 -538
rect 1687 -588 3287 -572
rect 3345 -538 4945 -500
rect 3345 -572 3361 -538
rect 4929 -572 4945 -538
rect 3345 -588 4945 -572
<< polycont >>
rect -4929 538 -3361 572
rect -3271 538 -1703 572
rect -1613 538 -45 572
rect 45 538 1613 572
rect 1703 538 3271 572
rect 3361 538 4929 572
rect -4929 -572 -3361 -538
rect -3271 -572 -1703 -538
rect -1613 -572 -45 -538
rect 45 -572 1613 -538
rect 1703 -572 3271 -538
rect 3361 -572 4929 -538
<< locali >>
rect -4945 538 -4929 572
rect -3361 538 -3345 572
rect -3287 538 -3271 572
rect -1703 538 -1687 572
rect -1629 538 -1613 572
rect -45 538 -29 572
rect 29 538 45 572
rect 1613 538 1629 572
rect 1687 538 1703 572
rect 3271 538 3287 572
rect 3345 538 3361 572
rect 4929 538 4945 572
rect -4991 488 -4957 504
rect -4991 -504 -4957 -488
rect -3333 488 -3299 504
rect -3333 -504 -3299 -488
rect -1675 488 -1641 504
rect -1675 -504 -1641 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 1641 488 1675 504
rect 1641 -504 1675 -488
rect 3299 488 3333 504
rect 3299 -504 3333 -488
rect 4957 488 4991 504
rect 4957 -504 4991 -488
rect -4945 -572 -4929 -538
rect -3361 -572 -3345 -538
rect -3287 -572 -3271 -538
rect -1703 -572 -1687 -538
rect -1629 -572 -1613 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 1613 -572 1629 -538
rect 1687 -572 1703 -538
rect 3271 -572 3287 -538
rect 3345 -572 3361 -538
rect 4929 -572 4945 -538
<< viali >>
rect -4929 538 -3361 572
rect -3271 538 -1703 572
rect -1613 538 -45 572
rect 45 538 1613 572
rect 1703 538 3271 572
rect 3361 538 4929 572
rect -4991 -488 -4957 488
rect -3333 -488 -3299 488
rect -1675 -488 -1641 488
rect -17 -488 17 488
rect 1641 -488 1675 488
rect 3299 -488 3333 488
rect 4957 -488 4991 488
rect -4929 -572 -3361 -538
rect -3271 -572 -1703 -538
rect -1613 -572 -45 -538
rect 45 -572 1613 -538
rect 1703 -572 3271 -538
rect 3361 -572 4929 -538
<< metal1 >>
rect -4941 572 -3349 578
rect -4941 538 -4929 572
rect -3361 538 -3349 572
rect -4941 532 -3349 538
rect -3283 572 -1691 578
rect -3283 538 -3271 572
rect -1703 538 -1691 572
rect -3283 532 -1691 538
rect -1625 572 -33 578
rect -1625 538 -1613 572
rect -45 538 -33 572
rect -1625 532 -33 538
rect 33 572 1625 578
rect 33 538 45 572
rect 1613 538 1625 572
rect 33 532 1625 538
rect 1691 572 3283 578
rect 1691 538 1703 572
rect 3271 538 3283 572
rect 1691 532 3283 538
rect 3349 572 4941 578
rect 3349 538 3361 572
rect 4929 538 4941 572
rect 3349 532 4941 538
rect -4997 488 -4951 500
rect -4997 -488 -4991 488
rect -4957 -488 -4951 488
rect -4997 -500 -4951 -488
rect -3339 488 -3293 500
rect -3339 -488 -3333 488
rect -3299 -488 -3293 488
rect -3339 -500 -3293 -488
rect -1681 488 -1635 500
rect -1681 -488 -1675 488
rect -1641 -488 -1635 488
rect -1681 -500 -1635 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 1635 488 1681 500
rect 1635 -488 1641 488
rect 1675 -488 1681 488
rect 1635 -500 1681 -488
rect 3293 488 3339 500
rect 3293 -488 3299 488
rect 3333 -488 3339 488
rect 3293 -500 3339 -488
rect 4951 488 4997 500
rect 4951 -488 4957 488
rect 4991 -488 4997 488
rect 4951 -500 4997 -488
rect -4941 -538 -3349 -532
rect -4941 -572 -4929 -538
rect -3361 -572 -3349 -538
rect -4941 -578 -3349 -572
rect -3283 -538 -1691 -532
rect -3283 -572 -3271 -538
rect -1703 -572 -1691 -538
rect -3283 -578 -1691 -572
rect -1625 -538 -33 -532
rect -1625 -572 -1613 -538
rect -45 -572 -33 -538
rect -1625 -578 -33 -572
rect 33 -538 1625 -532
rect 33 -572 45 -538
rect 1613 -572 1625 -538
rect 33 -578 1625 -572
rect 1691 -538 3283 -532
rect 1691 -572 1703 -538
rect 3271 -572 3283 -538
rect 1691 -578 3283 -572
rect 3349 -538 4941 -532
rect 3349 -572 3361 -538
rect 4929 -572 4941 -538
rect 3349 -578 4941 -572
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 8.0 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
