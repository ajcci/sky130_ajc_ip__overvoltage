magic
tech sky130A
timestamp 1712109191
<< pwell >>
rect -901 -379 901 379
<< mvnmos >>
rect -787 -250 -587 250
rect -558 -250 -358 250
rect -329 -250 -129 250
rect -100 -250 100 250
rect 129 -250 329 250
rect 358 -250 558 250
rect 587 -250 787 250
<< mvndiff >>
rect -816 244 -787 250
rect -816 -244 -810 244
rect -793 -244 -787 244
rect -816 -250 -787 -244
rect -587 244 -558 250
rect -587 -244 -581 244
rect -564 -244 -558 244
rect -587 -250 -558 -244
rect -358 244 -329 250
rect -358 -244 -352 244
rect -335 -244 -329 244
rect -358 -250 -329 -244
rect -129 244 -100 250
rect -129 -244 -123 244
rect -106 -244 -100 244
rect -129 -250 -100 -244
rect 100 244 129 250
rect 100 -244 106 244
rect 123 -244 129 244
rect 100 -250 129 -244
rect 329 244 358 250
rect 329 -244 335 244
rect 352 -244 358 244
rect 329 -250 358 -244
rect 558 244 587 250
rect 558 -244 564 244
rect 581 -244 587 244
rect 558 -250 587 -244
rect 787 244 816 250
rect 787 -244 793 244
rect 810 -244 816 244
rect 787 -250 816 -244
<< mvndiffc >>
rect -810 -244 -793 244
rect -581 -244 -564 244
rect -352 -244 -335 244
rect -123 -244 -106 244
rect 106 -244 123 244
rect 335 -244 352 244
rect 564 -244 581 244
rect 793 -244 810 244
<< mvpsubdiff >>
rect -883 355 883 361
rect -883 338 -829 355
rect 829 338 883 355
rect -883 332 883 338
rect -883 307 -854 332
rect -883 -307 -877 307
rect -860 -307 -854 307
rect 854 307 883 332
rect -883 -332 -854 -307
rect 854 -307 860 307
rect 877 -307 883 307
rect 854 -332 883 -307
rect -883 -338 883 -332
rect -883 -355 -829 -338
rect 829 -355 883 -338
rect -883 -361 883 -355
<< mvpsubdiffcont >>
rect -829 338 829 355
rect -877 -307 -860 307
rect 860 -307 877 307
rect -829 -355 829 -338
<< poly >>
rect -787 286 -587 294
rect -787 269 -779 286
rect -595 269 -587 286
rect -787 250 -587 269
rect -558 286 -358 294
rect -558 269 -550 286
rect -366 269 -358 286
rect -558 250 -358 269
rect -329 286 -129 294
rect -329 269 -321 286
rect -137 269 -129 286
rect -329 250 -129 269
rect -100 286 100 294
rect -100 269 -92 286
rect 92 269 100 286
rect -100 250 100 269
rect 129 286 329 294
rect 129 269 137 286
rect 321 269 329 286
rect 129 250 329 269
rect 358 286 558 294
rect 358 269 366 286
rect 550 269 558 286
rect 358 250 558 269
rect 587 286 787 294
rect 587 269 595 286
rect 779 269 787 286
rect 587 250 787 269
rect -787 -269 -587 -250
rect -787 -286 -779 -269
rect -595 -286 -587 -269
rect -787 -294 -587 -286
rect -558 -269 -358 -250
rect -558 -286 -550 -269
rect -366 -286 -358 -269
rect -558 -294 -358 -286
rect -329 -269 -129 -250
rect -329 -286 -321 -269
rect -137 -286 -129 -269
rect -329 -294 -129 -286
rect -100 -269 100 -250
rect -100 -286 -92 -269
rect 92 -286 100 -269
rect -100 -294 100 -286
rect 129 -269 329 -250
rect 129 -286 137 -269
rect 321 -286 329 -269
rect 129 -294 329 -286
rect 358 -269 558 -250
rect 358 -286 366 -269
rect 550 -286 558 -269
rect 358 -294 558 -286
rect 587 -269 787 -250
rect 587 -286 595 -269
rect 779 -286 787 -269
rect 587 -294 787 -286
<< polycont >>
rect -779 269 -595 286
rect -550 269 -366 286
rect -321 269 -137 286
rect -92 269 92 286
rect 137 269 321 286
rect 366 269 550 286
rect 595 269 779 286
rect -779 -286 -595 -269
rect -550 -286 -366 -269
rect -321 -286 -137 -269
rect -92 -286 92 -269
rect 137 -286 321 -269
rect 366 -286 550 -269
rect 595 -286 779 -269
<< locali >>
rect -877 338 -829 355
rect 829 338 877 355
rect -877 307 -860 338
rect 860 307 877 338
rect -787 269 -779 286
rect -595 269 -587 286
rect -558 269 -550 286
rect -366 269 -358 286
rect -329 269 -321 286
rect -137 269 -129 286
rect -100 269 -92 286
rect 92 269 100 286
rect 129 269 137 286
rect 321 269 329 286
rect 358 269 366 286
rect 550 269 558 286
rect 587 269 595 286
rect 779 269 787 286
rect -810 244 -793 252
rect -810 -252 -793 -244
rect -581 244 -564 252
rect -581 -252 -564 -244
rect -352 244 -335 252
rect -352 -252 -335 -244
rect -123 244 -106 252
rect -123 -252 -106 -244
rect 106 244 123 252
rect 106 -252 123 -244
rect 335 244 352 252
rect 335 -252 352 -244
rect 564 244 581 252
rect 564 -252 581 -244
rect 793 244 810 252
rect 793 -252 810 -244
rect -787 -286 -779 -269
rect -595 -286 -587 -269
rect -558 -286 -550 -269
rect -366 -286 -358 -269
rect -329 -286 -321 -269
rect -137 -286 -129 -269
rect -100 -286 -92 -269
rect 92 -286 100 -269
rect 129 -286 137 -269
rect 321 -286 329 -269
rect 358 -286 366 -269
rect 550 -286 558 -269
rect 587 -286 595 -269
rect 779 -286 787 -269
rect -877 -338 -860 -307
rect 860 -338 877 -307
rect -877 -355 -829 -338
rect 829 -355 877 -338
<< viali >>
rect -779 269 -595 286
rect -550 269 -366 286
rect -321 269 -137 286
rect -92 269 92 286
rect 137 269 321 286
rect 366 269 550 286
rect 595 269 779 286
rect -810 -244 -793 244
rect -581 -244 -564 244
rect -352 -244 -335 244
rect -123 -244 -106 244
rect 106 -244 123 244
rect 335 -244 352 244
rect 564 -244 581 244
rect 793 -244 810 244
rect -779 -286 -595 -269
rect -550 -286 -366 -269
rect -321 -286 -137 -269
rect -92 -286 92 -269
rect 137 -286 321 -269
rect 366 -286 550 -269
rect 595 -286 779 -269
<< metal1 >>
rect -785 286 -589 289
rect -785 269 -779 286
rect -595 269 -589 286
rect -785 266 -589 269
rect -556 286 -360 289
rect -556 269 -550 286
rect -366 269 -360 286
rect -556 266 -360 269
rect -327 286 -131 289
rect -327 269 -321 286
rect -137 269 -131 286
rect -327 266 -131 269
rect -98 286 98 289
rect -98 269 -92 286
rect 92 269 98 286
rect -98 266 98 269
rect 131 286 327 289
rect 131 269 137 286
rect 321 269 327 286
rect 131 266 327 269
rect 360 286 556 289
rect 360 269 366 286
rect 550 269 556 286
rect 360 266 556 269
rect 589 286 785 289
rect 589 269 595 286
rect 779 269 785 286
rect 589 266 785 269
rect -813 244 -790 250
rect -813 -244 -810 244
rect -793 -244 -790 244
rect -813 -250 -790 -244
rect -584 244 -561 250
rect -584 -244 -581 244
rect -564 -244 -561 244
rect -584 -250 -561 -244
rect -355 244 -332 250
rect -355 -244 -352 244
rect -335 -244 -332 244
rect -355 -250 -332 -244
rect -126 244 -103 250
rect -126 -244 -123 244
rect -106 -244 -103 244
rect -126 -250 -103 -244
rect 103 244 126 250
rect 103 -244 106 244
rect 123 -244 126 244
rect 103 -250 126 -244
rect 332 244 355 250
rect 332 -244 335 244
rect 352 -244 355 244
rect 332 -250 355 -244
rect 561 244 584 250
rect 561 -244 564 244
rect 581 -244 584 244
rect 561 -250 584 -244
rect 790 244 813 250
rect 790 -244 793 244
rect 810 -244 813 244
rect 790 -250 813 -244
rect -785 -269 -589 -266
rect -785 -286 -779 -269
rect -595 -286 -589 -269
rect -785 -289 -589 -286
rect -556 -269 -360 -266
rect -556 -286 -550 -269
rect -366 -286 -360 -269
rect -556 -289 -360 -286
rect -327 -269 -131 -266
rect -327 -286 -321 -269
rect -137 -286 -131 -269
rect -327 -289 -131 -286
rect -98 -269 98 -266
rect -98 -286 -92 -269
rect 92 -286 98 -269
rect -98 -289 98 -286
rect 131 -269 327 -266
rect 131 -286 137 -269
rect 321 -286 327 -269
rect 131 -289 327 -286
rect 360 -269 556 -266
rect 360 -286 366 -269
rect 550 -286 556 -269
rect 360 -289 556 -286
rect 589 -269 785 -266
rect 589 -286 595 -269
rect 779 -286 785 -269
rect 589 -289 785 -286
<< properties >>
string FIXED_BBOX -868 -346 868 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 2 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
