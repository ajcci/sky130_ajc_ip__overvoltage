magic
tech sky130A
timestamp 1712205713
<< pwell >>
rect -281 -155 281 155
<< nmos >>
rect -183 -50 -133 50
rect -104 -50 -54 50
rect -25 -50 25 50
rect 54 -50 104 50
rect 133 -50 183 50
<< ndiff >>
rect -212 44 -183 50
rect -212 -44 -206 44
rect -189 -44 -183 44
rect -212 -50 -183 -44
rect -133 44 -104 50
rect -133 -44 -127 44
rect -110 -44 -104 44
rect -133 -50 -104 -44
rect -54 44 -25 50
rect -54 -44 -48 44
rect -31 -44 -25 44
rect -54 -50 -25 -44
rect 25 44 54 50
rect 25 -44 31 44
rect 48 -44 54 44
rect 25 -50 54 -44
rect 104 44 133 50
rect 104 -44 110 44
rect 127 -44 133 44
rect 104 -50 133 -44
rect 183 44 212 50
rect 183 -44 189 44
rect 206 -44 212 44
rect 183 -50 212 -44
<< ndiffc >>
rect -206 -44 -189 44
rect -127 -44 -110 44
rect -48 -44 -31 44
rect 31 -44 48 44
rect 110 -44 127 44
rect 189 -44 206 44
<< psubdiff >>
rect -263 120 -215 137
rect 215 120 263 137
rect -263 89 -246 120
rect 246 89 263 120
rect -263 -120 -246 -89
rect 246 -120 263 -89
rect -263 -137 -215 -120
rect 215 -137 263 -120
<< psubdiffcont >>
rect -215 120 215 137
rect -263 -89 -246 89
rect 246 -89 263 89
rect -215 -137 215 -120
<< poly >>
rect -183 86 -133 94
rect -183 69 -175 86
rect -141 69 -133 86
rect -183 50 -133 69
rect -104 86 -54 94
rect -104 69 -96 86
rect -62 69 -54 86
rect -104 50 -54 69
rect -25 86 25 94
rect -25 69 -17 86
rect 17 69 25 86
rect -25 50 25 69
rect 54 86 104 94
rect 54 69 62 86
rect 96 69 104 86
rect 54 50 104 69
rect 133 86 183 94
rect 133 69 141 86
rect 175 69 183 86
rect 133 50 183 69
rect -183 -69 -133 -50
rect -183 -86 -175 -69
rect -141 -86 -133 -69
rect -183 -94 -133 -86
rect -104 -69 -54 -50
rect -104 -86 -96 -69
rect -62 -86 -54 -69
rect -104 -94 -54 -86
rect -25 -69 25 -50
rect -25 -86 -17 -69
rect 17 -86 25 -69
rect -25 -94 25 -86
rect 54 -69 104 -50
rect 54 -86 62 -69
rect 96 -86 104 -69
rect 54 -94 104 -86
rect 133 -69 183 -50
rect 133 -86 141 -69
rect 175 -86 183 -69
rect 133 -94 183 -86
<< polycont >>
rect -175 69 -141 86
rect -96 69 -62 86
rect -17 69 17 86
rect 62 69 96 86
rect 141 69 175 86
rect -175 -86 -141 -69
rect -96 -86 -62 -69
rect -17 -86 17 -69
rect 62 -86 96 -69
rect 141 -86 175 -69
<< locali >>
rect -263 120 -215 137
rect 215 120 263 137
rect -263 89 -246 120
rect 246 89 263 120
rect -183 69 -175 86
rect -141 69 -133 86
rect -104 69 -96 86
rect -62 69 -54 86
rect -25 69 -17 86
rect 17 69 25 86
rect 54 69 62 86
rect 96 69 104 86
rect 133 69 141 86
rect 175 69 183 86
rect -206 44 -189 52
rect -206 -52 -189 -44
rect -127 44 -110 52
rect -127 -52 -110 -44
rect -48 44 -31 52
rect -48 -52 -31 -44
rect 31 44 48 52
rect 31 -52 48 -44
rect 110 44 127 52
rect 110 -52 127 -44
rect 189 44 206 52
rect 189 -52 206 -44
rect -183 -86 -175 -69
rect -141 -86 -133 -69
rect -104 -86 -96 -69
rect -62 -86 -54 -69
rect -25 -86 -17 -69
rect 17 -86 25 -69
rect 54 -86 62 -69
rect 96 -86 104 -69
rect 133 -86 141 -69
rect 175 -86 183 -69
rect -263 -120 -246 -89
rect 246 -120 263 -89
rect -263 -137 -215 -120
rect 215 -137 263 -120
<< viali >>
rect -175 69 -141 86
rect -96 69 -62 86
rect -17 69 17 86
rect 62 69 96 86
rect 141 69 175 86
rect -206 -44 -189 44
rect -127 -44 -110 44
rect -48 -44 -31 44
rect 31 -44 48 44
rect 110 -44 127 44
rect 189 -44 206 44
rect -175 -86 -141 -69
rect -96 -86 -62 -69
rect -17 -86 17 -69
rect 62 -86 96 -69
rect 141 -86 175 -69
<< metal1 >>
rect -181 86 -135 89
rect -181 69 -175 86
rect -141 69 -135 86
rect -181 66 -135 69
rect -102 86 -56 89
rect -102 69 -96 86
rect -62 69 -56 86
rect -102 66 -56 69
rect -23 86 23 89
rect -23 69 -17 86
rect 17 69 23 86
rect -23 66 23 69
rect 56 86 102 89
rect 56 69 62 86
rect 96 69 102 86
rect 56 66 102 69
rect 135 86 181 89
rect 135 69 141 86
rect 175 69 181 86
rect 135 66 181 69
rect -209 44 -186 50
rect -209 -44 -206 44
rect -189 -44 -186 44
rect -209 -50 -186 -44
rect -130 44 -107 50
rect -130 -44 -127 44
rect -110 -44 -107 44
rect -130 -50 -107 -44
rect -51 44 -28 50
rect -51 -44 -48 44
rect -31 -44 -28 44
rect -51 -50 -28 -44
rect 28 44 51 50
rect 28 -44 31 44
rect 48 -44 51 44
rect 28 -50 51 -44
rect 107 44 130 50
rect 107 -44 110 44
rect 127 -44 130 44
rect 107 -50 130 -44
rect 186 44 209 50
rect 186 -44 189 44
rect 206 -44 209 44
rect 186 -50 209 -44
rect -181 -69 -135 -66
rect -181 -86 -175 -69
rect -141 -86 -135 -69
rect -181 -89 -135 -86
rect -102 -69 -56 -66
rect -102 -86 -96 -69
rect -62 -86 -56 -69
rect -102 -89 -56 -86
rect -23 -69 23 -66
rect -23 -86 -17 -69
rect 17 -86 23 -69
rect -23 -89 23 -86
rect 56 -69 102 -66
rect 56 -86 62 -69
rect 96 -86 102 -69
rect 56 -89 102 -86
rect 135 -69 181 -66
rect 135 -86 141 -69
rect 175 -86 181 -69
rect 135 -89 181 -86
<< properties >>
string FIXED_BBOX -254 -128 254 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.50 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
