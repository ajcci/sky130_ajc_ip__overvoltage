magic
tech sky130A
magscale 1 2
timestamp 1712338462
<< error_p >>
rect -4444 1342 -4370 1351
rect -4444 1286 -4435 1342
rect -4444 1277 -4370 1286
rect -4927 1094 -4853 1103
rect -4444 1094 -4370 1103
rect -4927 1038 -4918 1094
rect -4444 1038 -4435 1094
rect -4927 1029 -4853 1038
rect -4444 1029 -4370 1038
<< error_s >>
rect 3838 -7148 3861 -7147
rect 3838 -7196 3866 -7148
rect 7416 -7152 7480 -7151
rect 7411 -7179 7485 -7152
rect 7407 -7196 7489 -7179
rect 3829 -7201 3894 -7196
rect 3829 -7203 3843 -7201
rect 3856 -7203 3894 -7201
rect 7407 -7201 7480 -7196
rect 3829 -7205 3898 -7203
rect 3838 -7208 3898 -7205
rect 7407 -7207 7421 -7201
rect 3865 -7303 3866 -7208
rect 7411 -7212 7485 -7207
rect 9376 -7515 9381 -7460
rect 9376 -7520 9450 -7515
rect 9381 -7529 9386 -7520
rect 9376 -7584 9386 -7529
rect 9376 -7589 9450 -7584
<< locali >>
rect -4648 1400 -4520 1415
rect -4648 1302 -4633 1400
rect -4535 1302 -4520 1400
rect -4304 1400 -4240 1415
rect -4648 1287 -4520 1302
rect -4439 1331 -4375 1346
rect -4439 1297 -4424 1331
rect -4390 1297 -4375 1331
rect -4439 1282 -4375 1297
rect -4304 1302 -4289 1400
rect -4255 1302 -4240 1400
rect -4304 1287 -4240 1302
rect -3568 1284 -3510 1296
rect -3568 1250 -3556 1284
rect -3522 1250 -3510 1284
rect -3568 1238 -3510 1250
rect -3724 1142 -3596 1157
rect -3724 1044 -3709 1142
rect -3611 1044 -3596 1142
rect -3456 1142 -3392 1157
rect -3724 1029 -3596 1044
rect -3555 1078 -3491 1093
rect -3555 1044 -3540 1078
rect -3506 1044 -3491 1078
rect -3555 1029 -3491 1044
rect -3456 1044 -3441 1142
rect -3407 1044 -3392 1142
rect -3456 1029 -3392 1044
rect -3610 774 -3482 789
rect -3610 740 -3595 774
rect -3497 740 -3482 774
rect -3610 725 -3482 740
<< viali >>
rect -4633 1302 -4535 1400
rect -4424 1297 -4390 1331
rect -4289 1302 -4255 1400
rect -3556 1250 -3522 1284
rect -3709 1044 -3611 1142
rect -3540 1044 -3506 1078
rect -3441 1044 -3407 1142
rect -3595 740 -3497 774
<< metal1 >>
rect -4658 1414 -4510 1425
rect -4658 1288 -4647 1414
rect -4521 1288 -4510 1414
rect -4309 1414 -4235 1425
rect -4658 1277 -4510 1288
rect -4444 1340 -4370 1351
rect -4444 1288 -4433 1340
rect -4381 1288 -4370 1340
rect -4444 1277 -4370 1288
rect -4309 1288 -4298 1414
rect -4246 1288 -4235 1414
rect -4309 1277 -4235 1288
rect -3568 1284 -3510 1296
rect -3568 1250 -3556 1284
rect -3522 1250 -3510 1284
rect -3568 1238 -3510 1250
rect -4658 1166 -4510 1177
rect -4658 1040 -4647 1166
rect -4521 1040 -4510 1166
rect -4309 1166 -4235 1177
rect -4658 1029 -4510 1040
rect -4444 1092 -4370 1103
rect -4444 1040 -4433 1092
rect -4381 1040 -4370 1092
rect -4444 1029 -4370 1040
rect -4309 1040 -4298 1166
rect -4246 1040 -4235 1166
rect -4309 1029 -4235 1040
rect -4152 1151 -4024 1157
rect -4152 1035 -4146 1151
rect -4030 1035 -4024 1151
rect -3884 1151 -3820 1157
rect -4152 1029 -4024 1035
rect -3983 1087 -3919 1093
rect -3983 1035 -3977 1087
rect -3925 1035 -3919 1087
rect -3983 1029 -3919 1035
rect -3884 1035 -3878 1151
rect -3826 1035 -3820 1151
rect -3884 1029 -3820 1035
rect -3724 1151 -3596 1157
rect -3724 1035 -3718 1151
rect -3602 1035 -3596 1151
rect -3456 1151 -3392 1157
rect -3724 1029 -3596 1035
rect -3555 1087 -3491 1093
rect -3555 1035 -3549 1087
rect -3497 1035 -3491 1087
rect -3555 1029 -3491 1035
rect -3456 1035 -3450 1151
rect -3398 1035 -3392 1151
rect -3456 1029 -3392 1035
rect -3864 857 -3736 863
rect -3864 805 -3858 857
rect -3742 805 -3736 857
rect -3864 799 -3736 805
rect -3610 783 -3482 789
rect -4300 768 -4152 779
rect -4300 716 -4289 768
rect -4163 716 -4152 768
rect -3610 731 -3604 783
rect -3488 731 -3482 783
rect -3610 725 -3482 731
rect -4300 705 -4152 716
rect 3838 -3060 4648 -2912
rect 3838 -3874 4648 -3624
rect 3838 -4794 4648 -4438
rect 3838 -5608 4648 -5358
rect -27806 -10519 -27406 -10513
rect -27806 -10796 -27800 -10519
rect -27412 -10796 -27406 -10519
rect -27806 -10802 -27406 -10796
rect -19274 -10802 -10740 -10552
rect -28262 -10858 -27459 -10852
rect -28262 -11096 -28256 -10858
rect -27868 -11096 -27459 -10858
rect -28262 -11102 -27459 -11096
rect -19020 -11104 -10740 -10854
<< via1 >>
rect -4647 1400 -4521 1414
rect -4647 1302 -4633 1400
rect -4633 1302 -4535 1400
rect -4535 1302 -4521 1400
rect -4647 1288 -4521 1302
rect -4433 1331 -4381 1340
rect -4433 1297 -4424 1331
rect -4424 1297 -4390 1331
rect -4390 1297 -4381 1331
rect -4433 1288 -4381 1297
rect -4298 1400 -4246 1414
rect -4298 1302 -4289 1400
rect -4289 1302 -4255 1400
rect -4255 1302 -4246 1400
rect -4298 1288 -4246 1302
rect -4647 1040 -4521 1166
rect -4433 1040 -4381 1092
rect -4298 1040 -4246 1166
rect -4146 1035 -4030 1151
rect -3977 1035 -3925 1087
rect -3878 1035 -3826 1151
rect -3718 1142 -3602 1151
rect -3718 1044 -3709 1142
rect -3709 1044 -3611 1142
rect -3611 1044 -3602 1142
rect -3718 1035 -3602 1044
rect -3549 1078 -3497 1087
rect -3549 1044 -3540 1078
rect -3540 1044 -3506 1078
rect -3506 1044 -3497 1078
rect -3549 1035 -3497 1044
rect -3450 1142 -3398 1151
rect -3450 1044 -3441 1142
rect -3441 1044 -3407 1142
rect -3407 1044 -3398 1142
rect -3450 1035 -3398 1044
rect -3858 805 -3742 857
rect -4289 716 -4163 768
rect -3604 774 -3488 783
rect -3604 740 -3595 774
rect -3595 740 -3497 774
rect -3497 740 -3488 774
rect -3604 731 -3488 740
rect -27800 -10796 -27412 -10519
rect -28256 -11096 -27868 -10858
<< metal2 >>
rect -28262 10255 -27862 10398
rect -28262 10119 -27929 10255
rect -27868 10119 -27862 10255
rect -28262 -10858 -27862 10119
rect -27806 6812 -27406 10398
rect -19249 7756 -19185 7760
rect -19254 7751 -19180 7756
rect -19254 7687 -19249 7751
rect -19185 7687 -19180 7751
rect -27035 7147 -26979 7156
rect -27035 7082 -26979 7091
rect -27806 6676 -27478 6812
rect -27412 6676 -27406 6812
rect -27806 2314 -27406 6676
rect -27806 2178 -27478 2314
rect -27412 2178 -27406 2314
rect -27806 -10519 -27406 2178
rect -19254 607 -19180 7687
rect -17661 7151 -17597 7160
rect -18588 5514 -18528 5523
rect -18588 -8044 -18528 5454
rect -18293 5314 -18229 5323
rect -18293 2438 -18229 5250
rect -18293 2374 -18177 2438
rect -18241 -2878 -18177 2374
rect -17661 -2678 -17597 7087
rect -4658 1416 -4510 1425
rect -4658 1286 -4649 1416
rect -4519 1286 -4510 1416
rect -4309 1416 -4235 1425
rect -4658 1277 -4510 1286
rect -4444 1342 -4370 1351
rect -4444 1286 -4435 1342
rect -4379 1286 -4370 1342
rect -4444 1277 -4370 1286
rect -4309 1286 -4300 1416
rect -4244 1286 -4235 1416
rect -4309 1277 -4235 1286
rect -5142 1168 -4994 1177
rect -5142 1038 -5133 1168
rect -5003 1038 -4994 1168
rect -4793 1168 -4719 1177
rect -5142 1029 -4994 1038
rect -4927 1094 -4853 1103
rect -4927 1038 -4918 1094
rect -4862 1038 -4853 1094
rect -4927 1029 -4853 1038
rect -4793 1038 -4784 1168
rect -4728 1038 -4719 1168
rect -4793 1029 -4719 1038
rect -4658 1168 -4510 1177
rect -4658 1038 -4649 1168
rect -4519 1038 -4510 1168
rect -4309 1168 -4235 1177
rect -4658 1029 -4510 1038
rect -4444 1094 -4370 1103
rect -4444 1038 -4435 1094
rect -4379 1038 -4370 1094
rect -4444 1029 -4370 1038
rect -4309 1038 -4300 1168
rect -4244 1038 -4235 1168
rect -4309 1029 -4235 1038
rect -4152 1151 -4024 1157
rect -4152 1035 -4146 1151
rect -4030 1035 -4024 1151
rect -3884 1151 -3820 1157
rect -4152 1029 -4024 1035
rect -3983 1087 -3919 1093
rect -3983 1035 -3977 1087
rect -3925 1035 -3919 1087
rect -3983 1029 -3919 1035
rect -3884 1035 -3878 1151
rect -3826 1035 -3820 1151
rect -3884 1029 -3820 1035
rect -3724 1151 -3596 1157
rect -3724 1035 -3718 1151
rect -3602 1035 -3596 1151
rect -3456 1151 -3392 1157
rect -3724 1029 -3596 1035
rect -3555 1087 -3491 1093
rect -3555 1035 -3549 1087
rect -3497 1035 -3491 1087
rect -3555 1029 -3491 1035
rect -3456 1035 -3450 1151
rect -3398 1035 -3392 1151
rect -3456 1029 -3392 1035
rect -3864 857 -3736 863
rect -4784 814 -4636 823
rect -4784 758 -4775 814
rect -4645 758 -4636 814
rect -3864 805 -3858 857
rect -3742 805 -3736 857
rect -3864 799 -3736 805
rect -3610 783 -3482 789
rect -17531 605 -17457 753
rect -4784 749 -4636 758
rect -4300 770 -4152 779
rect -4300 714 -4291 770
rect -4161 714 -4152 770
rect -3610 731 -3604 783
rect -3488 731 -3482 783
rect -3610 725 -3482 731
rect -4300 705 -4152 714
rect -12959 -903 -12895 -894
rect -15351 -2196 -15287 -2068
rect -17666 -2734 -17657 -2678
rect -17601 -2734 -17592 -2678
rect -17661 -2738 -17597 -2734
rect -13162 -2745 -13084 -2709
rect -13162 -7524 -13098 -2745
rect -12959 -3378 -12895 -967
rect -12959 -3434 -12955 -3378
rect -12899 -3434 -12895 -3378
rect -12959 -3438 -12895 -3434
rect -12955 -3443 -12899 -3438
rect 3861 -7203 3865 -7196
rect 3838 -7368 3865 -7203
rect 7407 -7207 7416 -7196
rect 7480 -7207 7489 -7196
rect 3961 -7390 4025 -7248
rect -13162 -7580 -13158 -7524
rect -13102 -7580 -13098 -7524
rect -13162 -7584 -13098 -7580
rect 9381 -7520 9445 -7196
rect -13158 -7589 -13102 -7584
rect 9381 -7593 9445 -7584
rect -18588 -8100 -18586 -8044
rect -18530 -8100 -18528 -8044
rect -18588 -8102 -18528 -8100
rect -18586 -8109 -18530 -8102
rect -27806 -10796 -27800 -10519
rect -27412 -10796 -27406 -10519
rect -27806 -10802 -27406 -10796
rect -28262 -11096 -28256 -10858
rect -27868 -11096 -27862 -10858
rect -28262 -11102 -27862 -11096
<< via2 >>
rect -27929 10119 -27868 10255
rect -19249 7687 -19185 7751
rect -27035 7091 -26979 7147
rect -27478 6676 -27412 6812
rect -27478 2178 -27412 2314
rect -17661 7087 -17597 7151
rect -18588 5454 -18528 5514
rect -18293 5250 -18229 5314
rect -4649 1414 -4519 1416
rect -4649 1288 -4647 1414
rect -4647 1288 -4521 1414
rect -4521 1288 -4519 1414
rect -4649 1286 -4519 1288
rect -4435 1340 -4379 1342
rect -4435 1288 -4433 1340
rect -4433 1288 -4381 1340
rect -4381 1288 -4379 1340
rect -4435 1286 -4379 1288
rect -4300 1414 -4244 1416
rect -4300 1288 -4298 1414
rect -4298 1288 -4246 1414
rect -4246 1288 -4244 1414
rect -4300 1286 -4244 1288
rect -5133 1038 -5003 1168
rect -4918 1038 -4862 1094
rect -4784 1038 -4728 1168
rect -4649 1166 -4519 1168
rect -4649 1040 -4647 1166
rect -4647 1040 -4521 1166
rect -4521 1040 -4519 1166
rect -4649 1038 -4519 1040
rect -4435 1092 -4379 1094
rect -4435 1040 -4433 1092
rect -4433 1040 -4381 1092
rect -4381 1040 -4379 1092
rect -4435 1038 -4379 1040
rect -4300 1166 -4244 1168
rect -4300 1040 -4298 1166
rect -4298 1040 -4246 1166
rect -4246 1040 -4244 1166
rect -4300 1038 -4244 1040
rect -4775 758 -4645 814
rect -4291 768 -4161 770
rect -4291 716 -4289 768
rect -4289 716 -4163 768
rect -4163 716 -4161 768
rect -4291 714 -4161 716
rect -12959 -967 -12895 -903
rect -17657 -2734 -17601 -2678
rect -12955 -3434 -12899 -3378
rect 3838 -7203 3861 -7196
rect 7416 -7207 7480 -7196
rect -13158 -7580 -13102 -7524
rect 9381 -7584 9445 -7520
rect -18586 -8100 -18530 -8044
<< metal3 >>
rect -27935 10255 -27136 10261
rect -27935 10119 -27929 10255
rect -27868 10119 -27136 10255
rect -27935 10113 -27136 10119
rect -27218 7751 -19180 7756
rect -27218 7687 -19249 7751
rect -19185 7687 -19180 7751
rect -27218 7682 -19180 7687
rect -27040 7151 -26974 7152
rect -17666 7151 -17592 7156
rect -27040 7147 -17661 7151
rect -27040 7091 -27035 7147
rect -26979 7091 -17661 7147
rect -27040 7087 -17661 7091
rect -17597 7087 -17592 7151
rect -27040 7086 -26974 7087
rect -17666 7082 -17592 7087
rect -27484 6812 -27166 6818
rect -27484 6676 -27478 6812
rect -27412 6676 -27166 6812
rect -27484 6670 -27166 6676
rect -18593 5514 -18523 5519
rect -18593 5454 -18588 5514
rect -18528 5454 -18523 5514
rect -18593 5449 -18523 5454
rect -18298 5314 -18224 5319
rect -18298 5250 -18293 5314
rect -18229 5250 -18224 5314
rect -18298 5245 -18224 5250
rect -27484 2314 -26420 2320
rect -27484 2178 -27478 2314
rect -27412 2178 -26420 2314
rect -27484 2172 -26420 2178
rect -4658 1416 -4510 1425
rect -4658 1286 -4649 1416
rect -4519 1286 -4510 1416
rect -4309 1416 -4235 1425
rect -4658 1277 -4510 1286
rect -4444 1342 -4370 1351
rect -4444 1286 -4435 1342
rect -4379 1286 -4370 1342
rect -4444 1277 -4370 1286
rect -4309 1286 -4300 1416
rect -4244 1286 -4235 1416
rect -4309 1277 -4235 1286
rect -5142 1168 -4994 1177
rect -5142 1038 -5133 1168
rect -5003 1038 -4994 1168
rect -4793 1168 -4719 1177
rect -5142 1029 -4994 1038
rect -4927 1094 -4853 1103
rect -4927 1038 -4918 1094
rect -4862 1038 -4853 1094
rect -4927 1029 -4853 1038
rect -4793 1038 -4784 1168
rect -4728 1038 -4719 1168
rect -4793 1029 -4719 1038
rect -4658 1168 -4510 1177
rect -4658 1038 -4649 1168
rect -4519 1038 -4510 1168
rect -4309 1168 -4235 1177
rect -4658 1029 -4510 1038
rect -4444 1094 -4370 1103
rect -4444 1038 -4435 1094
rect -4379 1038 -4370 1094
rect -4444 1029 -4370 1038
rect -4309 1038 -4300 1168
rect -4244 1038 -4235 1168
rect -4309 1029 -4235 1038
rect -4784 814 -4636 823
rect -4784 758 -4775 814
rect -4645 758 -4636 814
rect -4784 749 -4636 758
rect -4300 770 -4152 779
rect -4300 714 -4291 770
rect -4161 714 -4152 770
rect -4300 705 -4152 714
rect -12964 -903 -12890 -898
rect -12964 -967 -12959 -903
rect -12895 -967 -12890 -903
rect -12964 -972 -12890 -967
rect -17662 -2674 -17596 -2673
rect -17662 -2678 -15348 -2674
rect -17662 -2734 -17657 -2678
rect -17601 -2734 -15348 -2678
rect -17662 -2738 -15348 -2734
rect -17662 -2739 -17596 -2738
rect -15414 -2793 -15348 -2738
rect -15414 -2858 -15412 -2793
rect -12960 -3374 -12894 -3373
rect -12960 -3378 -10740 -3374
rect -12960 -3434 -12955 -3378
rect -12899 -3434 -10740 -3378
rect -12960 -3438 -10740 -3434
rect -12960 -3439 -12894 -3438
rect 3838 -3750 4648 -3686
rect 3838 -7207 3861 -7203
rect 7480 -7207 7485 -7196
rect 3838 -7208 3866 -7207
rect 7411 -7212 7485 -7207
rect -13163 -7520 -13097 -7519
rect 9376 -7520 9450 -7515
rect -13163 -7524 -10740 -7520
rect -13163 -7580 -13158 -7524
rect -13102 -7580 -10740 -7524
rect -13163 -7584 -10740 -7580
rect 9445 -7584 9450 -7520
rect -13163 -7585 -13097 -7584
rect 9376 -7589 9450 -7584
rect -18591 -8042 -18525 -8039
rect -18591 -8044 -10740 -8042
rect -18591 -8100 -18586 -8044
rect -18530 -8100 -10740 -8044
rect -18591 -8102 -10740 -8100
rect -18591 -8105 -18525 -8102
use comparator  comparator_0
timestamp 1712334093
transform 1 0 -26517 0 1 2397
box -811 -518 11035 7864
use ibias_gen  ibias_gen_0
timestamp 1712334093
transform 1 0 -27321 0 1 -10450
box -138 -652 15828 11500
use rstring_mux  rstring_mux_0
timestamp 1712334093
transform 1 0 -16753 0 1 -15968
box -11632 -32 28451 9182
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 8 2112 0 1 1734
timestamp 1707688321
transform 1 0 -9540 0 1 -6297
box -66 -43 2178 1671
<< labels >>
flabel metal2 -17531 753 -17531 753 0 FreeSans 1200 0 0 0 itest
port 25 nsew
flabel metal2 s -18241 -2814 -18241 -2814 0 FreeSans 1200 0 0 0 vbg_1v2
port 26 nsew
flabel metal2 -15287 -2068 -15287 -2068 0 FreeSans 1200 0 0 0 ibg_200n
port 27 nsew
<< end >>
