magic
tech sky130A
magscale 1 2
timestamp 1712109191
<< pwell >>
rect -3898 -4082 3898 4082
<< psubdiff >>
rect -3862 4012 -3766 4046
rect 3766 4012 3862 4046
rect -3862 3950 -3828 4012
rect 3828 3950 3862 4012
rect -3862 -4012 -3828 -3950
rect 3828 -4012 3862 -3950
rect -3862 -4046 -3766 -4012
rect 3766 -4046 3862 -4012
<< psubdiffcont >>
rect -3766 4012 3766 4046
rect -3862 -3950 -3828 3950
rect 3828 -3950 3862 3950
rect -3766 -4046 3766 -4012
<< xpolycontact >>
rect -3732 3484 -3450 3916
rect -3732 -3916 -3450 -3484
rect -3354 3484 -3072 3916
rect -3354 -3916 -3072 -3484
rect -2976 3484 -2694 3916
rect -2976 -3916 -2694 -3484
rect -2598 3484 -2316 3916
rect -2598 -3916 -2316 -3484
rect -2220 3484 -1938 3916
rect -2220 -3916 -1938 -3484
rect -1842 3484 -1560 3916
rect -1842 -3916 -1560 -3484
rect -1464 3484 -1182 3916
rect -1464 -3916 -1182 -3484
rect -1086 3484 -804 3916
rect -1086 -3916 -804 -3484
rect -708 3484 -426 3916
rect -708 -3916 -426 -3484
rect -330 3484 -48 3916
rect -330 -3916 -48 -3484
rect 48 3484 330 3916
rect 48 -3916 330 -3484
rect 426 3484 708 3916
rect 426 -3916 708 -3484
rect 804 3484 1086 3916
rect 804 -3916 1086 -3484
rect 1182 3484 1464 3916
rect 1182 -3916 1464 -3484
rect 1560 3484 1842 3916
rect 1560 -3916 1842 -3484
rect 1938 3484 2220 3916
rect 1938 -3916 2220 -3484
rect 2316 3484 2598 3916
rect 2316 -3916 2598 -3484
rect 2694 3484 2976 3916
rect 2694 -3916 2976 -3484
rect 3072 3484 3354 3916
rect 3072 -3916 3354 -3484
rect 3450 3484 3732 3916
rect 3450 -3916 3732 -3484
<< xpolyres >>
rect -3732 -3484 -3450 3484
rect -3354 -3484 -3072 3484
rect -2976 -3484 -2694 3484
rect -2598 -3484 -2316 3484
rect -2220 -3484 -1938 3484
rect -1842 -3484 -1560 3484
rect -1464 -3484 -1182 3484
rect -1086 -3484 -804 3484
rect -708 -3484 -426 3484
rect -330 -3484 -48 3484
rect 48 -3484 330 3484
rect 426 -3484 708 3484
rect 804 -3484 1086 3484
rect 1182 -3484 1464 3484
rect 1560 -3484 1842 3484
rect 1938 -3484 2220 3484
rect 2316 -3484 2598 3484
rect 2694 -3484 2976 3484
rect 3072 -3484 3354 3484
rect 3450 -3484 3732 3484
<< locali >>
rect -3862 4012 -3766 4046
rect 3766 4012 3862 4046
rect -3862 3950 -3828 4012
rect 3828 3950 3862 4012
rect -3862 -4012 -3828 -3950
rect 3828 -4012 3862 -3950
rect -3862 -4046 -3766 -4012
rect 3766 -4046 3862 -4012
<< viali >>
rect -3716 3501 -3466 3898
rect -3338 3501 -3088 3898
rect -2960 3501 -2710 3898
rect -2582 3501 -2332 3898
rect -2204 3501 -1954 3898
rect -1826 3501 -1576 3898
rect -1448 3501 -1198 3898
rect -1070 3501 -820 3898
rect -692 3501 -442 3898
rect -314 3501 -64 3898
rect 64 3501 314 3898
rect 442 3501 692 3898
rect 820 3501 1070 3898
rect 1198 3501 1448 3898
rect 1576 3501 1826 3898
rect 1954 3501 2204 3898
rect 2332 3501 2582 3898
rect 2710 3501 2960 3898
rect 3088 3501 3338 3898
rect 3466 3501 3716 3898
rect -3716 -3898 -3466 -3501
rect -3338 -3898 -3088 -3501
rect -2960 -3898 -2710 -3501
rect -2582 -3898 -2332 -3501
rect -2204 -3898 -1954 -3501
rect -1826 -3898 -1576 -3501
rect -1448 -3898 -1198 -3501
rect -1070 -3898 -820 -3501
rect -692 -3898 -442 -3501
rect -314 -3898 -64 -3501
rect 64 -3898 314 -3501
rect 442 -3898 692 -3501
rect 820 -3898 1070 -3501
rect 1198 -3898 1448 -3501
rect 1576 -3898 1826 -3501
rect 1954 -3898 2204 -3501
rect 2332 -3898 2582 -3501
rect 2710 -3898 2960 -3501
rect 3088 -3898 3338 -3501
rect 3466 -3898 3716 -3501
<< metal1 >>
rect -3722 3898 -3460 3910
rect -3722 3501 -3716 3898
rect -3466 3501 -3460 3898
rect -3722 3489 -3460 3501
rect -3344 3898 -3082 3910
rect -3344 3501 -3338 3898
rect -3088 3501 -3082 3898
rect -3344 3489 -3082 3501
rect -2966 3898 -2704 3910
rect -2966 3501 -2960 3898
rect -2710 3501 -2704 3898
rect -2966 3489 -2704 3501
rect -2588 3898 -2326 3910
rect -2588 3501 -2582 3898
rect -2332 3501 -2326 3898
rect -2588 3489 -2326 3501
rect -2210 3898 -1948 3910
rect -2210 3501 -2204 3898
rect -1954 3501 -1948 3898
rect -2210 3489 -1948 3501
rect -1832 3898 -1570 3910
rect -1832 3501 -1826 3898
rect -1576 3501 -1570 3898
rect -1832 3489 -1570 3501
rect -1454 3898 -1192 3910
rect -1454 3501 -1448 3898
rect -1198 3501 -1192 3898
rect -1454 3489 -1192 3501
rect -1076 3898 -814 3910
rect -1076 3501 -1070 3898
rect -820 3501 -814 3898
rect -1076 3489 -814 3501
rect -698 3898 -436 3910
rect -698 3501 -692 3898
rect -442 3501 -436 3898
rect -698 3489 -436 3501
rect -320 3898 -58 3910
rect -320 3501 -314 3898
rect -64 3501 -58 3898
rect -320 3489 -58 3501
rect 58 3898 320 3910
rect 58 3501 64 3898
rect 314 3501 320 3898
rect 58 3489 320 3501
rect 436 3898 698 3910
rect 436 3501 442 3898
rect 692 3501 698 3898
rect 436 3489 698 3501
rect 814 3898 1076 3910
rect 814 3501 820 3898
rect 1070 3501 1076 3898
rect 814 3489 1076 3501
rect 1192 3898 1454 3910
rect 1192 3501 1198 3898
rect 1448 3501 1454 3898
rect 1192 3489 1454 3501
rect 1570 3898 1832 3910
rect 1570 3501 1576 3898
rect 1826 3501 1832 3898
rect 1570 3489 1832 3501
rect 1948 3898 2210 3910
rect 1948 3501 1954 3898
rect 2204 3501 2210 3898
rect 1948 3489 2210 3501
rect 2326 3898 2588 3910
rect 2326 3501 2332 3898
rect 2582 3501 2588 3898
rect 2326 3489 2588 3501
rect 2704 3898 2966 3910
rect 2704 3501 2710 3898
rect 2960 3501 2966 3898
rect 2704 3489 2966 3501
rect 3082 3898 3344 3910
rect 3082 3501 3088 3898
rect 3338 3501 3344 3898
rect 3082 3489 3344 3501
rect 3460 3898 3722 3910
rect 3460 3501 3466 3898
rect 3716 3501 3722 3898
rect 3460 3489 3722 3501
rect -3722 -3501 -3460 -3489
rect -3722 -3898 -3716 -3501
rect -3466 -3898 -3460 -3501
rect -3722 -3910 -3460 -3898
rect -3344 -3501 -3082 -3489
rect -3344 -3898 -3338 -3501
rect -3088 -3898 -3082 -3501
rect -3344 -3910 -3082 -3898
rect -2966 -3501 -2704 -3489
rect -2966 -3898 -2960 -3501
rect -2710 -3898 -2704 -3501
rect -2966 -3910 -2704 -3898
rect -2588 -3501 -2326 -3489
rect -2588 -3898 -2582 -3501
rect -2332 -3898 -2326 -3501
rect -2588 -3910 -2326 -3898
rect -2210 -3501 -1948 -3489
rect -2210 -3898 -2204 -3501
rect -1954 -3898 -1948 -3501
rect -2210 -3910 -1948 -3898
rect -1832 -3501 -1570 -3489
rect -1832 -3898 -1826 -3501
rect -1576 -3898 -1570 -3501
rect -1832 -3910 -1570 -3898
rect -1454 -3501 -1192 -3489
rect -1454 -3898 -1448 -3501
rect -1198 -3898 -1192 -3501
rect -1454 -3910 -1192 -3898
rect -1076 -3501 -814 -3489
rect -1076 -3898 -1070 -3501
rect -820 -3898 -814 -3501
rect -1076 -3910 -814 -3898
rect -698 -3501 -436 -3489
rect -698 -3898 -692 -3501
rect -442 -3898 -436 -3501
rect -698 -3910 -436 -3898
rect -320 -3501 -58 -3489
rect -320 -3898 -314 -3501
rect -64 -3898 -58 -3501
rect -320 -3910 -58 -3898
rect 58 -3501 320 -3489
rect 58 -3898 64 -3501
rect 314 -3898 320 -3501
rect 58 -3910 320 -3898
rect 436 -3501 698 -3489
rect 436 -3898 442 -3501
rect 692 -3898 698 -3501
rect 436 -3910 698 -3898
rect 814 -3501 1076 -3489
rect 814 -3898 820 -3501
rect 1070 -3898 1076 -3501
rect 814 -3910 1076 -3898
rect 1192 -3501 1454 -3489
rect 1192 -3898 1198 -3501
rect 1448 -3898 1454 -3501
rect 1192 -3910 1454 -3898
rect 1570 -3501 1832 -3489
rect 1570 -3898 1576 -3501
rect 1826 -3898 1832 -3501
rect 1570 -3910 1832 -3898
rect 1948 -3501 2210 -3489
rect 1948 -3898 1954 -3501
rect 2204 -3898 2210 -3501
rect 1948 -3910 2210 -3898
rect 2326 -3501 2588 -3489
rect 2326 -3898 2332 -3501
rect 2582 -3898 2588 -3501
rect 2326 -3910 2588 -3898
rect 2704 -3501 2966 -3489
rect 2704 -3898 2710 -3501
rect 2960 -3898 2966 -3501
rect 2704 -3910 2966 -3898
rect 3082 -3501 3344 -3489
rect 3082 -3898 3088 -3501
rect 3338 -3898 3344 -3501
rect 3082 -3910 3344 -3898
rect 3460 -3501 3722 -3489
rect 3460 -3898 3466 -3501
rect 3716 -3898 3722 -3501
rect 3460 -3910 3722 -3898
<< properties >>
string FIXED_BBOX -3845 -4029 3845 4029
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 35 m 1 nx 20 wmin 1.410 lmin 0.50 rho 2000 val 49.912k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
