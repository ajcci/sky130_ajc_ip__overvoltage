magic
tech sky130A
magscale 1 2
timestamp 1711690514
<< error_s >>
rect 18808 -2446 18826 -2432
rect 18826 -2466 18842 -2446
<< dnwell >>
rect 8363 -9837 36013 3064
<< nwell >>
rect 8283 2858 36093 3144
rect 8283 -9631 8569 2858
rect 35807 -9631 36093 2858
rect 8283 -9917 36093 -9631
<< pwell >>
rect 4522 -3169 6500 -1640
<< nsubdiff >>
rect 8320 3087 36056 3107
rect 8320 3053 8400 3087
rect 35976 3053 36056 3087
rect 8320 3033 36056 3053
rect 8320 3027 8394 3033
rect 8320 -9800 8340 3027
rect 8374 -9800 8394 3027
rect 8320 -9806 8394 -9800
rect 35982 3027 36056 3033
rect 35982 -9800 36002 3027
rect 36036 -9800 36056 3027
rect 35982 -9806 36056 -9800
rect 8320 -9826 36056 -9806
rect 8320 -9860 8400 -9826
rect 35976 -9860 36056 -9826
rect 8320 -9880 36056 -9860
<< mvpsubdiff >>
rect 5484 -2434 5665 -2401
rect 5484 -2468 5541 -2434
rect 5605 -2468 5665 -2434
rect 5484 -2492 5665 -2468
<< nsubdiffcont >>
rect 8400 3053 35976 3087
rect 8340 -9800 8374 3027
rect 36002 -9800 36036 3027
rect 8400 -9860 35976 -9826
<< mvpsubdiffcont >>
rect 5541 -2468 5605 -2434
<< locali >>
rect 8340 3053 8400 3087
rect 35976 3053 36036 3087
rect 8340 3027 8374 3053
rect 5516 -2434 5627 -2420
rect 5516 -2468 5541 -2434
rect 5605 -2468 5627 -2434
rect 5516 -2480 5627 -2468
rect 5547 -2520 5584 -2480
rect 36002 3027 36036 3053
rect 18706 -2478 18712 -2431
rect 8340 -9826 8374 -9800
rect 36002 -9826 36036 -9800
rect 8340 -9860 8400 -9826
rect 35976 -9860 36036 -9826
<< viali >>
rect 8340 -2485 8374 -2423
<< metal1 >>
rect 8329 -2423 8385 -2409
rect 8329 -2485 8340 -2423
rect 8374 -2485 8385 -2423
rect 8329 -2497 8385 -2485
rect 18545 -2609 18549 -2563
rect 18397 -2729 18443 -2725
rect 18555 -2729 18601 -2725
use flattenedmos  flattenedmos_0
timestamp 1711690227
transform 1 0 -1536 0 1 2458
box 19634 -5518 20560 -4674
<< labels >>
rlabel metal1 8329 -2444 8329 -2444 1 avdd
port 0 n
rlabel locali 5547 -2520 5547 -2520 1 avss
rlabel locali 18706 -2431 18706 -2431 7 vt
rlabel metal1 18549 -2563 18549 -2563 3 g
rlabel metal1 18397 -2729 18397 -2729 7 d
rlabel metal1 18601 -2729 18601 -2729 3 s
<< end >>
