magic
tech sky130A
magscale 1 2
timestamp 1712118495
<< nwell >>
rect -1603 -797 1603 797
<< mvpmos >>
rect -1345 -500 -945 500
rect -887 -500 -487 500
rect -429 -500 -29 500
rect 29 -500 429 500
rect 487 -500 887 500
rect 945 -500 1345 500
<< mvpdiff >>
rect -1403 488 -1345 500
rect -1403 -488 -1391 488
rect -1357 -488 -1345 488
rect -1403 -500 -1345 -488
rect -945 488 -887 500
rect -945 -488 -933 488
rect -899 -488 -887 488
rect -945 -500 -887 -488
rect -487 488 -429 500
rect -487 -488 -475 488
rect -441 -488 -429 488
rect -487 -500 -429 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 429 488 487 500
rect 429 -488 441 488
rect 475 -488 487 488
rect 429 -500 487 -488
rect 887 488 945 500
rect 887 -488 899 488
rect 933 -488 945 488
rect 887 -500 945 -488
rect 1345 488 1403 500
rect 1345 -488 1357 488
rect 1391 -488 1403 488
rect 1345 -500 1403 -488
<< mvpdiffc >>
rect -1391 -488 -1357 488
rect -933 -488 -899 488
rect -475 -488 -441 488
rect -17 -488 17 488
rect 441 -488 475 488
rect 899 -488 933 488
rect 1357 -488 1391 488
<< mvnsubdiff >>
rect -1537 719 1537 731
rect -1537 685 -1429 719
rect 1429 685 1537 719
rect -1537 673 1537 685
rect -1537 623 -1479 673
rect -1537 -623 -1525 623
rect -1491 -623 -1479 623
rect 1479 623 1537 673
rect -1537 -673 -1479 -623
rect 1479 -623 1491 623
rect 1525 -623 1537 623
rect 1479 -673 1537 -623
rect -1537 -685 1537 -673
rect -1537 -719 -1429 -685
rect 1429 -719 1537 -685
rect -1537 -731 1537 -719
<< mvnsubdiffcont >>
rect -1429 685 1429 719
rect -1525 -623 -1491 623
rect 1491 -623 1525 623
rect -1429 -719 1429 -685
<< poly >>
rect -1345 581 -945 597
rect -1345 547 -1329 581
rect -961 547 -945 581
rect -1345 500 -945 547
rect -887 581 -487 597
rect -887 547 -871 581
rect -503 547 -487 581
rect -887 500 -487 547
rect -429 581 -29 597
rect -429 547 -413 581
rect -45 547 -29 581
rect -429 500 -29 547
rect 29 581 429 597
rect 29 547 45 581
rect 413 547 429 581
rect 29 500 429 547
rect 487 581 887 597
rect 487 547 503 581
rect 871 547 887 581
rect 487 500 887 547
rect 945 581 1345 597
rect 945 547 961 581
rect 1329 547 1345 581
rect 945 500 1345 547
rect -1345 -547 -945 -500
rect -1345 -581 -1329 -547
rect -961 -581 -945 -547
rect -1345 -597 -945 -581
rect -887 -547 -487 -500
rect -887 -581 -871 -547
rect -503 -581 -487 -547
rect -887 -597 -487 -581
rect -429 -547 -29 -500
rect -429 -581 -413 -547
rect -45 -581 -29 -547
rect -429 -597 -29 -581
rect 29 -547 429 -500
rect 29 -581 45 -547
rect 413 -581 429 -547
rect 29 -597 429 -581
rect 487 -547 887 -500
rect 487 -581 503 -547
rect 871 -581 887 -547
rect 487 -597 887 -581
rect 945 -547 1345 -500
rect 945 -581 961 -547
rect 1329 -581 1345 -547
rect 945 -597 1345 -581
<< polycont >>
rect -1329 547 -961 581
rect -871 547 -503 581
rect -413 547 -45 581
rect 45 547 413 581
rect 503 547 871 581
rect 961 547 1329 581
rect -1329 -581 -961 -547
rect -871 -581 -503 -547
rect -413 -581 -45 -547
rect 45 -581 413 -547
rect 503 -581 871 -547
rect 961 -581 1329 -547
<< locali >>
rect -1525 685 -1429 719
rect 1429 685 1525 719
rect -1525 623 -1491 685
rect 1491 623 1525 685
rect -1345 547 -1329 581
rect -961 547 -945 581
rect -887 547 -871 581
rect -503 547 -487 581
rect -429 547 -413 581
rect -45 547 -29 581
rect 29 547 45 581
rect 413 547 429 581
rect 487 547 503 581
rect 871 547 887 581
rect 945 547 961 581
rect 1329 547 1345 581
rect -1391 488 -1357 504
rect -1391 -504 -1357 -488
rect -933 488 -899 504
rect -933 -504 -899 -488
rect -475 488 -441 504
rect -475 -504 -441 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 441 488 475 504
rect 441 -504 475 -488
rect 899 488 933 504
rect 899 -504 933 -488
rect 1357 488 1391 504
rect 1357 -504 1391 -488
rect -1345 -581 -1329 -547
rect -961 -581 -945 -547
rect -887 -581 -871 -547
rect -503 -581 -487 -547
rect -429 -581 -413 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 413 -581 429 -547
rect 487 -581 503 -547
rect 871 -581 887 -547
rect 945 -581 961 -547
rect 1329 -581 1345 -547
rect -1525 -685 -1491 -623
rect 1491 -685 1525 -623
rect -1525 -719 -1429 -685
rect 1429 -719 1525 -685
<< viali >>
rect -1329 547 -961 581
rect -871 547 -503 581
rect -413 547 -45 581
rect 45 547 413 581
rect 503 547 871 581
rect 961 547 1329 581
rect -1391 -488 -1357 488
rect -933 -488 -899 488
rect -475 -488 -441 488
rect -17 -488 17 488
rect 441 -488 475 488
rect 899 -488 933 488
rect 1357 -488 1391 488
rect -1329 -581 -961 -547
rect -871 -581 -503 -547
rect -413 -581 -45 -547
rect 45 -581 413 -547
rect 503 -581 871 -547
rect 961 -581 1329 -547
<< metal1 >>
rect -1341 581 -949 587
rect -1341 547 -1329 581
rect -961 547 -949 581
rect -1341 541 -949 547
rect -883 581 -491 587
rect -883 547 -871 581
rect -503 547 -491 581
rect -883 541 -491 547
rect -425 581 -33 587
rect -425 547 -413 581
rect -45 547 -33 581
rect -425 541 -33 547
rect 33 581 425 587
rect 33 547 45 581
rect 413 547 425 581
rect 33 541 425 547
rect 491 581 883 587
rect 491 547 503 581
rect 871 547 883 581
rect 491 541 883 547
rect 949 581 1341 587
rect 949 547 961 581
rect 1329 547 1341 581
rect 949 541 1341 547
rect -1397 488 -1351 500
rect -1397 -488 -1391 488
rect -1357 -488 -1351 488
rect -1397 -500 -1351 -488
rect -939 488 -893 500
rect -939 -488 -933 488
rect -899 -488 -893 488
rect -939 -500 -893 -488
rect -481 488 -435 500
rect -481 -488 -475 488
rect -441 -488 -435 488
rect -481 -500 -435 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 435 488 481 500
rect 435 -488 441 488
rect 475 -488 481 488
rect 435 -500 481 -488
rect 893 488 939 500
rect 893 -488 899 488
rect 933 -488 939 488
rect 893 -500 939 -488
rect 1351 488 1397 500
rect 1351 -488 1357 488
rect 1391 -488 1397 488
rect 1351 -500 1397 -488
rect -1341 -547 -949 -541
rect -1341 -581 -1329 -547
rect -961 -581 -949 -547
rect -1341 -587 -949 -581
rect -883 -547 -491 -541
rect -883 -581 -871 -547
rect -503 -581 -491 -547
rect -883 -587 -491 -581
rect -425 -547 -33 -541
rect -425 -581 -413 -547
rect -45 -581 -33 -547
rect -425 -587 -33 -581
rect 33 -547 425 -541
rect 33 -581 45 -547
rect 413 -581 425 -547
rect 33 -587 425 -581
rect 491 -547 883 -541
rect 491 -581 503 -547
rect 871 -581 883 -547
rect 491 -587 883 -581
rect 949 -547 1341 -541
rect 949 -581 961 -547
rect 1329 -581 1341 -547
rect 949 -587 1341 -581
<< properties >>
string FIXED_BBOX -1508 -702 1508 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 2 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
