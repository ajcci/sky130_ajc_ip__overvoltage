magic
tech sky130A
timestamp 1711636687
<< nwell >>
rect -5088 -214 5088 214
<< mvpmos >>
rect -4959 23 -4159 65
rect -4130 23 -3330 65
rect -3301 23 -2501 65
rect -2472 23 -1672 65
rect -1643 23 -843 65
rect -814 23 -14 65
rect 14 23 814 65
rect 843 23 1643 65
rect 1672 23 2472 65
rect 2501 23 3301 65
rect 3330 23 4130 65
rect 4159 23 4959 65
rect -4959 -101 -4159 -59
rect -4130 -101 -3330 -59
rect -3301 -101 -2501 -59
rect -2472 -101 -1672 -59
rect -1643 -101 -843 -59
rect -814 -101 -14 -59
rect 14 -101 814 -59
rect 843 -101 1643 -59
rect 1672 -101 2472 -59
rect 2501 -101 3301 -59
rect 3330 -101 4130 -59
rect 4159 -101 4959 -59
<< mvpdiff >>
rect -4988 59 -4959 65
rect -4988 29 -4982 59
rect -4965 29 -4959 59
rect -4988 23 -4959 29
rect -4159 59 -4130 65
rect -4159 29 -4153 59
rect -4136 29 -4130 59
rect -4159 23 -4130 29
rect -3330 59 -3301 65
rect -3330 29 -3324 59
rect -3307 29 -3301 59
rect -3330 23 -3301 29
rect -2501 59 -2472 65
rect -2501 29 -2495 59
rect -2478 29 -2472 59
rect -2501 23 -2472 29
rect -1672 59 -1643 65
rect -1672 29 -1666 59
rect -1649 29 -1643 59
rect -1672 23 -1643 29
rect -843 59 -814 65
rect -843 29 -837 59
rect -820 29 -814 59
rect -843 23 -814 29
rect -14 59 14 65
rect -14 29 -8 59
rect 8 29 14 59
rect -14 23 14 29
rect 814 59 843 65
rect 814 29 820 59
rect 837 29 843 59
rect 814 23 843 29
rect 1643 59 1672 65
rect 1643 29 1649 59
rect 1666 29 1672 59
rect 1643 23 1672 29
rect 2472 59 2501 65
rect 2472 29 2478 59
rect 2495 29 2501 59
rect 2472 23 2501 29
rect 3301 59 3330 65
rect 3301 29 3307 59
rect 3324 29 3330 59
rect 3301 23 3330 29
rect 4130 59 4159 65
rect 4130 29 4136 59
rect 4153 29 4159 59
rect 4130 23 4159 29
rect 4959 59 4988 65
rect 4959 29 4965 59
rect 4982 29 4988 59
rect 4959 23 4988 29
rect -4988 -65 -4959 -59
rect -4988 -95 -4982 -65
rect -4965 -95 -4959 -65
rect -4988 -101 -4959 -95
rect -4159 -65 -4130 -59
rect -4159 -95 -4153 -65
rect -4136 -95 -4130 -65
rect -4159 -101 -4130 -95
rect -3330 -65 -3301 -59
rect -3330 -95 -3324 -65
rect -3307 -95 -3301 -65
rect -3330 -101 -3301 -95
rect -2501 -65 -2472 -59
rect -2501 -95 -2495 -65
rect -2478 -95 -2472 -65
rect -2501 -101 -2472 -95
rect -1672 -65 -1643 -59
rect -1672 -95 -1666 -65
rect -1649 -95 -1643 -65
rect -1672 -101 -1643 -95
rect -843 -65 -814 -59
rect -843 -95 -837 -65
rect -820 -95 -814 -65
rect -843 -101 -814 -95
rect -14 -65 14 -59
rect -14 -95 -8 -65
rect 8 -95 14 -65
rect -14 -101 14 -95
rect 814 -65 843 -59
rect 814 -95 820 -65
rect 837 -95 843 -65
rect 814 -101 843 -95
rect 1643 -65 1672 -59
rect 1643 -95 1649 -65
rect 1666 -95 1672 -65
rect 1643 -101 1672 -95
rect 2472 -65 2501 -59
rect 2472 -95 2478 -65
rect 2495 -95 2501 -65
rect 2472 -101 2501 -95
rect 3301 -65 3330 -59
rect 3301 -95 3307 -65
rect 3324 -95 3330 -65
rect 3301 -101 3330 -95
rect 4130 -65 4159 -59
rect 4130 -95 4136 -65
rect 4153 -95 4159 -65
rect 4130 -101 4159 -95
rect 4959 -65 4988 -59
rect 4959 -95 4965 -65
rect 4982 -95 4988 -65
rect 4959 -101 4988 -95
<< mvpdiffc >>
rect -4982 29 -4965 59
rect -4153 29 -4136 59
rect -3324 29 -3307 59
rect -2495 29 -2478 59
rect -1666 29 -1649 59
rect -837 29 -820 59
rect -8 29 8 59
rect 820 29 837 59
rect 1649 29 1666 59
rect 2478 29 2495 59
rect 3307 29 3324 59
rect 4136 29 4153 59
rect 4965 29 4982 59
rect -4982 -95 -4965 -65
rect -4153 -95 -4136 -65
rect -3324 -95 -3307 -65
rect -2495 -95 -2478 -65
rect -1666 -95 -1649 -65
rect -837 -95 -820 -65
rect -8 -95 8 -65
rect 820 -95 837 -65
rect 1649 -95 1666 -65
rect 2478 -95 2495 -65
rect 3307 -95 3324 -65
rect 4136 -95 4153 -65
rect 4965 -95 4982 -65
<< mvnsubdiff >>
rect -5055 175 5055 181
rect -5055 158 -5001 175
rect 5001 158 5055 175
rect -5055 152 5055 158
rect -5055 127 -5026 152
rect -5055 -127 -5049 127
rect -5032 -127 -5026 127
rect 5026 127 5055 152
rect -5055 -152 -5026 -127
rect 5026 -127 5032 127
rect 5049 -127 5055 127
rect 5026 -152 5055 -127
rect -5055 -158 5055 -152
rect -5055 -175 -5001 -158
rect 5001 -175 5055 -158
rect -5055 -181 5055 -175
<< mvnsubdiffcont >>
rect -5001 158 5001 175
rect -5049 -127 -5032 127
rect 5032 -127 5049 127
rect -5001 -175 5001 -158
<< poly >>
rect -4959 106 -4159 114
rect -4959 89 -4951 106
rect -4167 89 -4159 106
rect -4959 65 -4159 89
rect -4130 106 -3330 114
rect -4130 89 -4122 106
rect -3338 89 -3330 106
rect -4130 65 -3330 89
rect -3301 106 -2501 114
rect -3301 89 -3293 106
rect -2509 89 -2501 106
rect -3301 65 -2501 89
rect -2472 106 -1672 114
rect -2472 89 -2464 106
rect -1680 89 -1672 106
rect -2472 65 -1672 89
rect -1643 106 -843 114
rect -1643 89 -1635 106
rect -851 89 -843 106
rect -1643 65 -843 89
rect -814 106 -14 114
rect -814 89 -806 106
rect -22 89 -14 106
rect -814 65 -14 89
rect 14 106 814 114
rect 14 89 22 106
rect 806 89 814 106
rect 14 65 814 89
rect 843 106 1643 114
rect 843 89 851 106
rect 1635 89 1643 106
rect 843 65 1643 89
rect 1672 106 2472 114
rect 1672 89 1680 106
rect 2464 89 2472 106
rect 1672 65 2472 89
rect 2501 106 3301 114
rect 2501 89 2509 106
rect 3293 89 3301 106
rect 2501 65 3301 89
rect 3330 106 4130 114
rect 3330 89 3338 106
rect 4122 89 4130 106
rect 3330 65 4130 89
rect 4159 106 4959 114
rect 4159 89 4167 106
rect 4951 89 4959 106
rect 4159 65 4959 89
rect -4959 10 -4159 23
rect -4130 10 -3330 23
rect -3301 10 -2501 23
rect -2472 10 -1672 23
rect -1643 10 -843 23
rect -814 10 -14 23
rect 14 10 814 23
rect 843 10 1643 23
rect 1672 10 2472 23
rect 2501 10 3301 23
rect 3330 10 4130 23
rect 4159 10 4959 23
rect -4959 -18 -4159 -10
rect -4959 -35 -4951 -18
rect -4167 -35 -4159 -18
rect -4959 -59 -4159 -35
rect -4130 -18 -3330 -10
rect -4130 -35 -4122 -18
rect -3338 -35 -3330 -18
rect -4130 -59 -3330 -35
rect -3301 -18 -2501 -10
rect -3301 -35 -3293 -18
rect -2509 -35 -2501 -18
rect -3301 -59 -2501 -35
rect -2472 -18 -1672 -10
rect -2472 -35 -2464 -18
rect -1680 -35 -1672 -18
rect -2472 -59 -1672 -35
rect -1643 -18 -843 -10
rect -1643 -35 -1635 -18
rect -851 -35 -843 -18
rect -1643 -59 -843 -35
rect -814 -18 -14 -10
rect -814 -35 -806 -18
rect -22 -35 -14 -18
rect -814 -59 -14 -35
rect 14 -18 814 -10
rect 14 -35 22 -18
rect 806 -35 814 -18
rect 14 -59 814 -35
rect 843 -18 1643 -10
rect 843 -35 851 -18
rect 1635 -35 1643 -18
rect 843 -59 1643 -35
rect 1672 -18 2472 -10
rect 1672 -35 1680 -18
rect 2464 -35 2472 -18
rect 1672 -59 2472 -35
rect 2501 -18 3301 -10
rect 2501 -35 2509 -18
rect 3293 -35 3301 -18
rect 2501 -59 3301 -35
rect 3330 -18 4130 -10
rect 3330 -35 3338 -18
rect 4122 -35 4130 -18
rect 3330 -59 4130 -35
rect 4159 -18 4959 -10
rect 4159 -35 4167 -18
rect 4951 -35 4959 -18
rect 4159 -59 4959 -35
rect -4959 -114 -4159 -101
rect -4130 -114 -3330 -101
rect -3301 -114 -2501 -101
rect -2472 -114 -1672 -101
rect -1643 -114 -843 -101
rect -814 -114 -14 -101
rect 14 -114 814 -101
rect 843 -114 1643 -101
rect 1672 -114 2472 -101
rect 2501 -114 3301 -101
rect 3330 -114 4130 -101
rect 4159 -114 4959 -101
<< polycont >>
rect -4951 89 -4167 106
rect -4122 89 -3338 106
rect -3293 89 -2509 106
rect -2464 89 -1680 106
rect -1635 89 -851 106
rect -806 89 -22 106
rect 22 89 806 106
rect 851 89 1635 106
rect 1680 89 2464 106
rect 2509 89 3293 106
rect 3338 89 4122 106
rect 4167 89 4951 106
rect -4951 -35 -4167 -18
rect -4122 -35 -3338 -18
rect -3293 -35 -2509 -18
rect -2464 -35 -1680 -18
rect -1635 -35 -851 -18
rect -806 -35 -22 -18
rect 22 -35 806 -18
rect 851 -35 1635 -18
rect 1680 -35 2464 -18
rect 2509 -35 3293 -18
rect 3338 -35 4122 -18
rect 4167 -35 4951 -18
<< locali >>
rect -5049 158 -5001 175
rect 5001 158 5049 175
rect -5049 127 -5032 158
rect 5032 127 5049 158
rect -4959 89 -4951 106
rect -4167 89 -4159 106
rect -4130 89 -4122 106
rect -3338 89 -3330 106
rect -3301 89 -3293 106
rect -2509 89 -2501 106
rect -2472 89 -2464 106
rect -1680 89 -1672 106
rect -1643 89 -1635 106
rect -851 89 -843 106
rect -814 89 -806 106
rect -22 89 -14 106
rect 14 89 22 106
rect 806 89 814 106
rect 843 89 851 106
rect 1635 89 1643 106
rect 1672 89 1680 106
rect 2464 89 2472 106
rect 2501 89 2509 106
rect 3293 89 3301 106
rect 3330 89 3338 106
rect 4122 89 4130 106
rect 4159 89 4167 106
rect 4951 89 4959 106
rect -4982 59 -4965 67
rect -4982 21 -4965 29
rect -4153 59 -4136 67
rect -4153 21 -4136 29
rect -3324 59 -3307 67
rect -3324 21 -3307 29
rect -2495 59 -2478 67
rect -2495 21 -2478 29
rect -1666 59 -1649 67
rect -1666 21 -1649 29
rect -837 59 -820 67
rect -837 21 -820 29
rect -8 59 8 67
rect -8 21 8 29
rect 820 59 837 67
rect 820 21 837 29
rect 1649 59 1666 67
rect 1649 21 1666 29
rect 2478 59 2495 67
rect 2478 21 2495 29
rect 3307 59 3324 67
rect 3307 21 3324 29
rect 4136 59 4153 67
rect 4136 21 4153 29
rect 4965 59 4982 67
rect 4965 21 4982 29
rect -4959 -35 -4951 -18
rect -4167 -35 -4159 -18
rect -4130 -35 -4122 -18
rect -3338 -35 -3330 -18
rect -3301 -35 -3293 -18
rect -2509 -35 -2501 -18
rect -2472 -35 -2464 -18
rect -1680 -35 -1672 -18
rect -1643 -35 -1635 -18
rect -851 -35 -843 -18
rect -814 -35 -806 -18
rect -22 -35 -14 -18
rect 14 -35 22 -18
rect 806 -35 814 -18
rect 843 -35 851 -18
rect 1635 -35 1643 -18
rect 1672 -35 1680 -18
rect 2464 -35 2472 -18
rect 2501 -35 2509 -18
rect 3293 -35 3301 -18
rect 3330 -35 3338 -18
rect 4122 -35 4130 -18
rect 4159 -35 4167 -18
rect 4951 -35 4959 -18
rect -4982 -65 -4965 -57
rect -4982 -103 -4965 -95
rect -4153 -65 -4136 -57
rect -4153 -103 -4136 -95
rect -3324 -65 -3307 -57
rect -3324 -103 -3307 -95
rect -2495 -65 -2478 -57
rect -2495 -103 -2478 -95
rect -1666 -65 -1649 -57
rect -1666 -103 -1649 -95
rect -837 -65 -820 -57
rect -837 -103 -820 -95
rect -8 -65 8 -57
rect -8 -103 8 -95
rect 820 -65 837 -57
rect 820 -103 837 -95
rect 1649 -65 1666 -57
rect 1649 -103 1666 -95
rect 2478 -65 2495 -57
rect 2478 -103 2495 -95
rect 3307 -65 3324 -57
rect 3307 -103 3324 -95
rect 4136 -65 4153 -57
rect 4136 -103 4153 -95
rect 4965 -65 4982 -57
rect 4965 -103 4982 -95
rect -5049 -158 -5032 -127
rect 5032 -158 5049 -127
rect -5049 -175 -5001 -158
rect 5001 -175 5049 -158
<< viali >>
rect -4951 89 -4167 106
rect -4122 89 -3338 106
rect -3293 89 -2509 106
rect -2464 89 -1680 106
rect -1635 89 -851 106
rect -806 89 -22 106
rect 22 89 806 106
rect 851 89 1635 106
rect 1680 89 2464 106
rect 2509 89 3293 106
rect 3338 89 4122 106
rect 4167 89 4951 106
rect -4982 29 -4965 59
rect -4153 29 -4136 59
rect -3324 29 -3307 59
rect -2495 29 -2478 59
rect -1666 29 -1649 59
rect -837 29 -820 59
rect -8 29 8 59
rect 820 29 837 59
rect 1649 29 1666 59
rect 2478 29 2495 59
rect 3307 29 3324 59
rect 4136 29 4153 59
rect 4965 29 4982 59
rect -4951 -35 -4167 -18
rect -4122 -35 -3338 -18
rect -3293 -35 -2509 -18
rect -2464 -35 -1680 -18
rect -1635 -35 -851 -18
rect -806 -35 -22 -18
rect 22 -35 806 -18
rect 851 -35 1635 -18
rect 1680 -35 2464 -18
rect 2509 -35 3293 -18
rect 3338 -35 4122 -18
rect 4167 -35 4951 -18
rect -4982 -95 -4965 -65
rect -4153 -95 -4136 -65
rect -3324 -95 -3307 -65
rect -2495 -95 -2478 -65
rect -1666 -95 -1649 -65
rect -837 -95 -820 -65
rect -8 -95 8 -65
rect 820 -95 837 -65
rect 1649 -95 1666 -65
rect 2478 -95 2495 -65
rect 3307 -95 3324 -65
rect 4136 -95 4153 -65
rect 4965 -95 4982 -65
<< metal1 >>
rect -4957 106 -4161 109
rect -4957 89 -4951 106
rect -4167 89 -4161 106
rect -4957 86 -4161 89
rect -4128 106 -3332 109
rect -4128 89 -4122 106
rect -3338 89 -3332 106
rect -4128 86 -3332 89
rect -3299 106 -2503 109
rect -3299 89 -3293 106
rect -2509 89 -2503 106
rect -3299 86 -2503 89
rect -2470 106 -1674 109
rect -2470 89 -2464 106
rect -1680 89 -1674 106
rect -2470 86 -1674 89
rect -1641 106 -845 109
rect -1641 89 -1635 106
rect -851 89 -845 106
rect -1641 86 -845 89
rect -812 106 -16 109
rect -812 89 -806 106
rect -22 89 -16 106
rect -812 86 -16 89
rect 16 106 812 109
rect 16 89 22 106
rect 806 89 812 106
rect 16 86 812 89
rect 845 106 1641 109
rect 845 89 851 106
rect 1635 89 1641 106
rect 845 86 1641 89
rect 1674 106 2470 109
rect 1674 89 1680 106
rect 2464 89 2470 106
rect 1674 86 2470 89
rect 2503 106 3299 109
rect 2503 89 2509 106
rect 3293 89 3299 106
rect 2503 86 3299 89
rect 3332 106 4128 109
rect 3332 89 3338 106
rect 4122 89 4128 106
rect 3332 86 4128 89
rect 4161 106 4957 109
rect 4161 89 4167 106
rect 4951 89 4957 106
rect 4161 86 4957 89
rect -4985 59 -4962 65
rect -4985 29 -4982 59
rect -4965 29 -4962 59
rect -4985 23 -4962 29
rect -4156 59 -4133 65
rect -4156 29 -4153 59
rect -4136 29 -4133 59
rect -4156 23 -4133 29
rect -3327 59 -3304 65
rect -3327 29 -3324 59
rect -3307 29 -3304 59
rect -3327 23 -3304 29
rect -2498 59 -2475 65
rect -2498 29 -2495 59
rect -2478 29 -2475 59
rect -2498 23 -2475 29
rect -1669 59 -1646 65
rect -1669 29 -1666 59
rect -1649 29 -1646 59
rect -1669 23 -1646 29
rect -840 59 -817 65
rect -840 29 -837 59
rect -820 29 -817 59
rect -840 23 -817 29
rect -11 59 11 65
rect -11 29 -8 59
rect 8 29 11 59
rect -11 23 11 29
rect 817 59 840 65
rect 817 29 820 59
rect 837 29 840 59
rect 817 23 840 29
rect 1646 59 1669 65
rect 1646 29 1649 59
rect 1666 29 1669 59
rect 1646 23 1669 29
rect 2475 59 2498 65
rect 2475 29 2478 59
rect 2495 29 2498 59
rect 2475 23 2498 29
rect 3304 59 3327 65
rect 3304 29 3307 59
rect 3324 29 3327 59
rect 3304 23 3327 29
rect 4133 59 4156 65
rect 4133 29 4136 59
rect 4153 29 4156 59
rect 4133 23 4156 29
rect 4962 59 4985 65
rect 4962 29 4965 59
rect 4982 29 4985 59
rect 4962 23 4985 29
rect -4957 -18 -4161 -15
rect -4957 -35 -4951 -18
rect -4167 -35 -4161 -18
rect -4957 -38 -4161 -35
rect -4128 -18 -3332 -15
rect -4128 -35 -4122 -18
rect -3338 -35 -3332 -18
rect -4128 -38 -3332 -35
rect -3299 -18 -2503 -15
rect -3299 -35 -3293 -18
rect -2509 -35 -2503 -18
rect -3299 -38 -2503 -35
rect -2470 -18 -1674 -15
rect -2470 -35 -2464 -18
rect -1680 -35 -1674 -18
rect -2470 -38 -1674 -35
rect -1641 -18 -845 -15
rect -1641 -35 -1635 -18
rect -851 -35 -845 -18
rect -1641 -38 -845 -35
rect -812 -18 -16 -15
rect -812 -35 -806 -18
rect -22 -35 -16 -18
rect -812 -38 -16 -35
rect 16 -18 812 -15
rect 16 -35 22 -18
rect 806 -35 812 -18
rect 16 -38 812 -35
rect 845 -18 1641 -15
rect 845 -35 851 -18
rect 1635 -35 1641 -18
rect 845 -38 1641 -35
rect 1674 -18 2470 -15
rect 1674 -35 1680 -18
rect 2464 -35 2470 -18
rect 1674 -38 2470 -35
rect 2503 -18 3299 -15
rect 2503 -35 2509 -18
rect 3293 -35 3299 -18
rect 2503 -38 3299 -35
rect 3332 -18 4128 -15
rect 3332 -35 3338 -18
rect 4122 -35 4128 -18
rect 3332 -38 4128 -35
rect 4161 -18 4957 -15
rect 4161 -35 4167 -18
rect 4951 -35 4957 -18
rect 4161 -38 4957 -35
rect -4985 -65 -4962 -59
rect -4985 -95 -4982 -65
rect -4965 -95 -4962 -65
rect -4985 -101 -4962 -95
rect -4156 -65 -4133 -59
rect -4156 -95 -4153 -65
rect -4136 -95 -4133 -65
rect -4156 -101 -4133 -95
rect -3327 -65 -3304 -59
rect -3327 -95 -3324 -65
rect -3307 -95 -3304 -65
rect -3327 -101 -3304 -95
rect -2498 -65 -2475 -59
rect -2498 -95 -2495 -65
rect -2478 -95 -2475 -65
rect -2498 -101 -2475 -95
rect -1669 -65 -1646 -59
rect -1669 -95 -1666 -65
rect -1649 -95 -1646 -65
rect -1669 -101 -1646 -95
rect -840 -65 -817 -59
rect -840 -95 -837 -65
rect -820 -95 -817 -65
rect -840 -101 -817 -95
rect -11 -65 11 -59
rect -11 -95 -8 -65
rect 8 -95 11 -65
rect -11 -101 11 -95
rect 817 -65 840 -59
rect 817 -95 820 -65
rect 837 -95 840 -65
rect 817 -101 840 -95
rect 1646 -65 1669 -59
rect 1646 -95 1649 -65
rect 1666 -95 1669 -65
rect 1646 -101 1669 -95
rect 2475 -65 2498 -59
rect 2475 -95 2478 -65
rect 2495 -95 2498 -65
rect 2475 -101 2498 -95
rect 3304 -65 3327 -59
rect 3304 -95 3307 -65
rect 3324 -95 3327 -65
rect 3304 -101 3327 -95
rect 4133 -65 4156 -59
rect 4133 -95 4136 -65
rect 4153 -95 4156 -65
rect 4133 -101 4156 -95
rect 4962 -65 4985 -59
rect 4962 -95 4965 -65
rect 4982 -95 4985 -65
rect 4962 -101 4985 -95
<< properties >>
string FIXED_BBOX -5041 -166 5041 166
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 8.0 m 2 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
