magic
tech sky130A
magscale 1 2
timestamp 1711636687
<< pwell >>
rect -377 -308 377 308
<< mvnmos >>
rect -149 -50 -29 50
rect 29 -50 149 50
<< mvndiff >>
rect -207 38 -149 50
rect -207 -38 -195 38
rect -161 -38 -149 38
rect -207 -50 -149 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 149 38 207 50
rect 149 -38 161 38
rect 195 -38 207 38
rect 149 -50 207 -38
<< mvndiffc >>
rect -195 -38 -161 38
rect -17 -38 17 38
rect 161 -38 195 38
<< mvpsubdiff >>
rect -341 260 341 272
rect -341 226 -233 260
rect 233 226 341 260
rect -341 214 341 226
rect -341 164 -283 214
rect -341 -164 -329 164
rect -295 -164 -283 164
rect 283 164 341 214
rect -341 -214 -283 -164
rect 283 -164 295 164
rect 329 -164 341 164
rect 283 -214 341 -164
rect -341 -226 341 -214
rect -341 -260 -233 -226
rect 233 -260 341 -226
rect -341 -272 341 -260
<< mvpsubdiffcont >>
rect -233 226 233 260
rect -329 -164 -295 164
rect 295 -164 329 164
rect -233 -260 233 -226
<< poly >>
rect -149 122 -29 138
rect -149 88 -133 122
rect -45 88 -29 122
rect -149 50 -29 88
rect 29 122 149 138
rect 29 88 45 122
rect 133 88 149 122
rect 29 50 149 88
rect -149 -88 -29 -50
rect -149 -122 -133 -88
rect -45 -122 -29 -88
rect -149 -138 -29 -122
rect 29 -88 149 -50
rect 29 -122 45 -88
rect 133 -122 149 -88
rect 29 -138 149 -122
<< polycont >>
rect -133 88 -45 122
rect 45 88 133 122
rect -133 -122 -45 -88
rect 45 -122 133 -88
<< locali >>
rect -329 226 -233 260
rect 233 226 329 260
rect -329 164 -295 226
rect 295 164 329 226
rect -149 88 -133 122
rect -45 88 -29 122
rect 29 88 45 122
rect 133 88 149 122
rect -195 38 -161 54
rect -195 -54 -161 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 161 38 195 54
rect 161 -54 195 -38
rect -149 -122 -133 -88
rect -45 -122 -29 -88
rect 29 -122 45 -88
rect 133 -122 149 -88
rect -329 -226 -295 -164
rect 295 -226 329 -164
rect -329 -260 -233 -226
rect 233 -260 329 -226
<< viali >>
rect -133 88 -45 122
rect 45 88 133 122
rect -195 -38 -161 38
rect -17 -38 17 38
rect 161 -38 195 38
rect -133 -122 -45 -88
rect 45 -122 133 -88
<< metal1 >>
rect -145 122 -33 128
rect -145 88 -133 122
rect -45 88 -33 122
rect -145 82 -33 88
rect 33 122 145 128
rect 33 88 45 122
rect 133 88 145 122
rect 33 82 145 88
rect -201 38 -155 50
rect -201 -38 -195 38
rect -161 -38 -155 38
rect -201 -50 -155 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 155 38 201 50
rect 155 -38 161 38
rect 195 -38 201 38
rect 155 -50 201 -38
rect -145 -88 -33 -82
rect -145 -122 -133 -88
rect -45 -122 -33 -88
rect -145 -128 -33 -122
rect 33 -88 145 -82
rect 33 -122 45 -88
rect 133 -122 145 -88
rect 33 -128 145 -122
<< properties >>
string FIXED_BBOX -312 -243 312 243
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 0.6 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
