magic
tech sky130A
magscale 1 2
timestamp 1712369776
<< metal3 >>
rect -3186 18812 3186 18840
rect -3186 12788 3102 18812
rect 3166 12788 3186 18812
rect -3186 12760 3186 12788
rect -3186 12492 3186 12520
rect -3186 6468 3102 12492
rect 3166 6468 3186 12492
rect -3186 6440 3186 6468
rect -3186 6172 3186 6200
rect -3186 148 3102 6172
rect 3166 148 3186 6172
rect -3186 120 3186 148
rect -3186 -148 3186 -120
rect -3186 -6172 3102 -148
rect 3166 -6172 3186 -148
rect -3186 -6200 3186 -6172
rect -3186 -6468 3186 -6440
rect -3186 -12492 3102 -6468
rect 3166 -12492 3186 -6468
rect -3186 -12520 3186 -12492
rect -3186 -12788 3186 -12760
rect -3186 -18812 3102 -12788
rect 3166 -18812 3186 -12788
rect -3186 -18840 3186 -18812
<< via3 >>
rect 3102 12788 3166 18812
rect 3102 6468 3166 12492
rect 3102 148 3166 6172
rect 3102 -6172 3166 -148
rect 3102 -12492 3166 -6468
rect 3102 -18812 3166 -12788
<< mimcap >>
rect -3146 18760 2854 18800
rect -3146 12840 -3106 18760
rect 2814 12840 2854 18760
rect -3146 12800 2854 12840
rect -3146 12440 2854 12480
rect -3146 6520 -3106 12440
rect 2814 6520 2854 12440
rect -3146 6480 2854 6520
rect -3146 6120 2854 6160
rect -3146 200 -3106 6120
rect 2814 200 2854 6120
rect -3146 160 2854 200
rect -3146 -200 2854 -160
rect -3146 -6120 -3106 -200
rect 2814 -6120 2854 -200
rect -3146 -6160 2854 -6120
rect -3146 -6520 2854 -6480
rect -3146 -12440 -3106 -6520
rect 2814 -12440 2854 -6520
rect -3146 -12480 2854 -12440
rect -3146 -12840 2854 -12800
rect -3146 -18760 -3106 -12840
rect 2814 -18760 2854 -12840
rect -3146 -18800 2854 -18760
<< mimcapcontact >>
rect -3106 12840 2814 18760
rect -3106 6520 2814 12440
rect -3106 200 2814 6120
rect -3106 -6120 2814 -200
rect -3106 -12440 2814 -6520
rect -3106 -18760 2814 -12840
<< metal4 >>
rect -198 18761 -94 18960
rect 3082 18812 3186 18960
rect -3107 18760 2815 18761
rect -3107 12840 -3106 18760
rect 2814 12840 2815 18760
rect -3107 12839 2815 12840
rect -198 12441 -94 12839
rect 3082 12788 3102 18812
rect 3166 12788 3186 18812
rect 3082 12492 3186 12788
rect -3107 12440 2815 12441
rect -3107 6520 -3106 12440
rect 2814 6520 2815 12440
rect -3107 6519 2815 6520
rect -198 6121 -94 6519
rect 3082 6468 3102 12492
rect 3166 6468 3186 12492
rect 3082 6172 3186 6468
rect -3107 6120 2815 6121
rect -3107 200 -3106 6120
rect 2814 200 2815 6120
rect -3107 199 2815 200
rect -198 -199 -94 199
rect 3082 148 3102 6172
rect 3166 148 3186 6172
rect 3082 -148 3186 148
rect -3107 -200 2815 -199
rect -3107 -6120 -3106 -200
rect 2814 -6120 2815 -200
rect -3107 -6121 2815 -6120
rect -198 -6519 -94 -6121
rect 3082 -6172 3102 -148
rect 3166 -6172 3186 -148
rect 3082 -6468 3186 -6172
rect -3107 -6520 2815 -6519
rect -3107 -12440 -3106 -6520
rect 2814 -12440 2815 -6520
rect -3107 -12441 2815 -12440
rect -198 -12839 -94 -12441
rect 3082 -12492 3102 -6468
rect 3166 -12492 3186 -6468
rect 3082 -12788 3186 -12492
rect -3107 -12840 2815 -12839
rect -3107 -18760 -3106 -12840
rect 2814 -18760 2815 -12840
rect -3107 -18761 2815 -18760
rect -198 -18960 -94 -18761
rect 3082 -18812 3102 -12788
rect 3166 -18812 3186 -12788
rect 3082 -18960 3186 -18812
<< properties >>
string FIXED_BBOX -3186 12760 2894 18840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
