magic
tech sky130A
magscale 1 2
timestamp 1712450145
<< nwell >>
rect 53 1015 99 1082
<< pwell >>
rect 622 374 714 425
rect 92 29 138 96
rect 408 29 454 96
rect 724 29 770 96
<< viali >>
rect 41 1093 2165 1127
rect 41 631 2165 665
rect 80 436 940 470
rect 80 -16 940 18
<< metal1 >>
rect -66 1127 2272 1138
rect -66 1093 41 1127
rect 2165 1093 2272 1127
rect -66 1082 2272 1093
rect -66 676 -10 1082
rect 53 1015 99 1082
rect 369 1015 415 1082
rect 685 1015 731 1082
rect 1001 1015 1047 1082
rect 1317 1015 1363 1082
rect 1633 1015 1679 1082
rect 1949 1015 1995 1082
rect 202 980 266 986
rect 202 876 208 980
rect 260 876 266 980
rect 202 870 266 876
rect 518 980 582 986
rect 518 876 524 980
rect 576 876 582 980
rect 518 870 582 876
rect 834 980 898 986
rect 834 876 840 980
rect 892 876 898 980
rect 834 870 898 876
rect 1150 980 1214 986
rect 1150 876 1156 980
rect 1208 876 1214 980
rect 1150 870 1214 876
rect 1466 980 1530 986
rect 1466 876 1472 980
rect 1524 876 1530 980
rect 1466 870 1530 876
rect 1782 980 1846 986
rect 1782 876 1788 980
rect 1840 876 1846 980
rect 1782 870 1846 876
rect 2098 980 2162 986
rect 2098 876 2104 980
rect 2156 876 2162 980
rect 2098 870 2162 876
rect 325 776 389 782
rect 325 774 331 776
rect 201 728 331 774
rect 325 724 331 728
rect 383 774 389 776
rect 1177 776 1241 782
rect 1177 774 1183 776
rect 383 728 899 774
rect 1149 728 1183 774
rect 383 724 389 728
rect 325 718 389 724
rect 1177 724 1183 728
rect 1235 774 1241 776
rect 1846 774 1910 779
rect 1235 728 1373 774
rect 1781 773 2005 774
rect 1781 728 1852 773
rect 1235 724 1241 728
rect 1177 718 1241 724
rect 1531 676 1623 728
rect 1846 721 1852 728
rect 1904 728 2005 773
rect 1904 721 1910 728
rect 1846 715 1910 721
rect 2216 676 2272 1082
rect -66 665 2272 676
rect -66 631 41 665
rect 2165 631 2272 665
rect -66 620 2272 631
rect -27 470 1047 481
rect -27 436 80 470
rect 940 436 1047 470
rect -27 425 1047 436
rect -27 29 29 425
rect 330 386 394 392
rect 240 328 306 374
rect 330 334 336 386
rect 388 334 394 386
rect 330 328 394 334
rect 484 384 548 390
rect 484 332 490 384
rect 542 332 548 384
rect 622 374 714 425
rect 803 386 867 392
rect 484 326 548 332
rect 803 334 809 386
rect 861 334 867 386
rect 803 328 867 334
rect 241 262 305 268
rect 241 210 247 262
rect 299 210 305 262
rect 241 204 305 210
rect 557 262 621 268
rect 557 210 563 262
rect 615 210 621 262
rect 557 204 621 210
rect 873 262 937 268
rect 873 210 879 262
rect 931 210 937 262
rect 873 204 937 210
rect 92 29 138 96
rect 408 29 454 96
rect 724 29 770 96
rect 991 29 1047 425
rect -27 18 1047 29
rect -27 -16 80 18
rect 940 -16 1047 18
rect -27 -27 1047 -16
<< via1 >>
rect 208 876 260 980
rect 524 876 576 980
rect 840 876 892 980
rect 1156 876 1208 980
rect 1472 876 1524 980
rect 1788 876 1840 980
rect 2104 876 2156 980
rect 331 724 383 776
rect 1183 724 1235 776
rect 1852 721 1904 773
rect 336 334 388 386
rect 490 332 542 384
rect 809 334 861 386
rect 247 210 299 262
rect 563 210 615 262
rect 879 210 931 262
<< metal2 >>
rect 197 981 271 990
rect 197 875 206 981
rect 262 875 271 981
rect 197 866 271 875
rect 513 981 587 990
rect 513 875 522 981
rect 578 875 587 981
rect 513 866 587 875
rect 829 981 903 990
rect 829 875 838 981
rect 894 875 903 981
rect 1145 981 1219 990
rect 1145 929 1154 981
rect 829 866 903 875
rect 1043 875 1154 929
rect 1210 875 1219 981
rect 1043 869 1219 875
rect 215 268 271 866
rect 325 776 389 782
rect 325 724 331 776
rect 383 724 389 776
rect 325 718 389 724
rect 333 392 389 718
rect 619 714 679 723
rect 1043 712 1103 869
rect 1145 866 1219 869
rect 1461 981 1535 990
rect 1461 875 1470 981
rect 1526 875 1535 981
rect 1777 981 1851 990
rect 1645 926 1701 933
rect 1461 866 1535 875
rect 1643 924 1703 926
rect 1643 868 1645 924
rect 1701 868 1703 924
rect 1043 656 1045 712
rect 1101 656 1103 712
rect 1043 654 1103 656
rect 1177 776 1241 782
rect 1177 724 1183 776
rect 1235 724 1241 776
rect 1177 718 1241 724
rect 619 645 679 654
rect 1045 647 1101 654
rect 481 565 559 574
rect 481 505 490 565
rect 550 505 559 565
rect 481 496 559 505
rect 330 386 394 392
rect 492 390 548 496
rect 330 334 336 386
rect 388 334 394 386
rect 330 328 394 334
rect 484 384 548 390
rect 621 394 677 645
rect 1177 563 1237 718
rect 1177 507 1179 563
rect 1235 507 1237 563
rect 798 394 872 397
rect 621 388 872 394
rect 621 387 807 388
rect 484 332 490 384
rect 542 332 548 384
rect 484 326 548 332
rect 591 332 807 387
rect 863 332 872 388
rect 591 331 872 332
rect 591 268 647 331
rect 798 323 872 331
rect 215 265 305 268
rect 557 265 647 268
rect 215 262 647 265
rect 215 234 247 262
rect 241 210 247 234
rect 299 210 563 262
rect 615 230 647 262
rect 873 262 937 268
rect 873 256 879 262
rect 931 256 937 262
rect 615 210 621 230
rect 241 209 621 210
rect 241 204 305 209
rect 557 204 621 209
rect 873 204 878 256
rect 934 204 937 256
rect 1177 255 1237 507
rect 878 191 934 200
rect 1177 186 1237 195
rect 1643 258 1703 868
rect 1777 875 1786 981
rect 1842 875 1851 981
rect 1777 866 1851 875
rect 2093 981 2167 990
rect 2093 875 2102 981
rect 2158 875 2167 981
rect 2093 866 2167 875
rect 1846 773 1910 779
rect 1846 721 1852 773
rect 1904 721 1910 773
rect 1846 715 1910 721
rect 1848 388 1908 715
rect 1848 332 1850 388
rect 1906 332 1908 388
rect 1848 330 1908 332
rect 1850 323 1906 330
rect 1643 189 1703 198
<< via2 >>
rect 206 980 262 981
rect 206 876 208 980
rect 208 876 260 980
rect 260 876 262 980
rect 206 875 262 876
rect 522 980 578 981
rect 522 876 524 980
rect 524 876 576 980
rect 576 876 578 980
rect 522 875 578 876
rect 838 980 894 981
rect 838 876 840 980
rect 840 876 892 980
rect 892 876 894 980
rect 838 875 894 876
rect 1154 980 1210 981
rect 1154 876 1156 980
rect 1156 876 1208 980
rect 1208 876 1210 980
rect 1154 875 1210 876
rect 619 654 679 714
rect 1470 980 1526 981
rect 1470 876 1472 980
rect 1472 876 1524 980
rect 1524 876 1526 980
rect 1470 875 1526 876
rect 1645 868 1701 924
rect 1045 656 1101 712
rect 490 505 550 565
rect 1179 507 1235 563
rect 807 386 863 388
rect 807 334 809 386
rect 809 334 861 386
rect 861 334 863 386
rect 807 332 863 334
rect 878 210 879 256
rect 879 210 931 256
rect 931 210 934 256
rect 878 200 934 210
rect 1177 195 1237 255
rect 1786 980 1842 981
rect 1786 876 1788 980
rect 1788 876 1840 980
rect 1840 876 1842 980
rect 1786 875 1842 876
rect 2102 980 2158 981
rect 2102 876 2104 980
rect 2104 876 2156 980
rect 2156 876 2158 980
rect 2102 875 2158 876
rect 1850 332 1906 388
rect 1643 198 1703 258
<< metal3 >>
rect 197 981 271 990
rect 197 875 206 981
rect 262 926 271 981
rect 513 981 587 990
rect 513 926 522 981
rect 262 875 522 926
rect 578 926 587 981
rect 829 981 903 990
rect 829 926 838 981
rect 578 875 838 926
rect 894 875 903 981
rect 197 866 903 875
rect 1145 981 1219 990
rect 1145 875 1154 981
rect 1210 926 1219 981
rect 1461 981 1535 990
rect 1461 926 1470 981
rect 1210 875 1470 926
rect 1526 875 1535 981
rect 1777 981 1851 990
rect 1145 866 1535 875
rect 1640 926 1706 929
rect 1777 926 1786 981
rect 1640 924 1786 926
rect 1640 868 1645 924
rect 1701 875 1786 924
rect 1842 926 1851 981
rect 2093 981 2167 990
rect 2093 926 2102 981
rect 1842 875 2102 926
rect 2158 875 2167 981
rect 1701 868 2167 875
rect 1640 866 2167 868
rect 1640 863 1706 866
rect 614 714 684 719
rect 1040 714 1106 717
rect 614 654 619 714
rect 679 712 1106 714
rect 679 656 1045 712
rect 1101 656 1106 712
rect 679 654 1106 656
rect 614 649 684 654
rect 1040 651 1106 654
rect 485 565 555 570
rect 1174 565 1240 568
rect 485 505 490 565
rect 550 563 1240 565
rect 550 507 1179 563
rect 1235 507 1240 563
rect 550 505 1240 507
rect 485 500 555 505
rect 1174 502 1240 505
rect 798 390 872 397
rect 1845 390 1911 393
rect 798 388 1911 390
rect 798 332 807 388
rect 863 332 1850 388
rect 1906 332 1911 388
rect 798 330 1911 332
rect 798 323 872 330
rect 1845 327 1911 330
rect 873 258 939 261
rect 1172 258 1242 260
rect 1638 258 1708 263
rect 873 256 1643 258
rect 873 200 878 256
rect 934 255 1643 256
rect 934 200 1177 255
rect 873 198 1177 200
rect 873 195 939 198
rect 1172 195 1177 198
rect 1237 198 1643 255
rect 1703 198 1708 258
rect 1237 195 1242 198
rect 1172 190 1242 195
rect 1638 193 1708 198
use sky130_fd_pr__nfet_01v8_SCV3UK  sky130_fd_pr__nfet_01v8_SCV3UK_1
timestamp 1712422266
transform 1 0 510 0 1 227
box -562 -279 562 279
use sky130_fd_pr__pfet_01v8_BZXTE7  sky130_fd_pr__pfet_01v8_BZXTE7_0
timestamp 1712422266
transform 1 0 1103 0 1 879
box -1194 -284 1194 284
<< labels >>
flabel metal1 -27 481 -27 481 0 FreeSans 800 0 0 0 dvss
port 4 nsew
flabel metal1 -66 1138 -66 1138 0 FreeSans 800 0 0 0 dvdd
port 1 nsew
flabel metal2 333 548 333 548 0 FreeSans 800 0 0 0 in
port 2 nsew
flabel metal2 1703 534 1703 534 0 FreeSans 800 0 0 0 out
port 3 nsew
flabel metal2 215 546 215 546 0 FreeSans 800 0 0 0 m
<< end >>
