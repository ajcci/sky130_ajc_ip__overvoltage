magic
tech sky130A
magscale 1 2
timestamp 1711823137
<< error_s >>
rect -1039 6252 -965 6261
rect -1039 6196 -1030 6252
rect -1039 6187 -965 6196
<< locali >>
rect 102 7501 166 7516
rect 102 7467 117 7501
rect 151 7467 166 7501
rect 102 7452 166 7467
rect 1760 7501 1824 7516
rect 1760 7467 1775 7501
rect 1809 7467 1824 7501
rect 1760 7452 1824 7467
rect 5076 7501 5140 7516
rect 5076 7467 5091 7501
rect 5125 7467 5140 7501
rect 5076 7452 5140 7467
rect 8392 7501 8456 7516
rect 8392 7467 8407 7501
rect 8441 7467 8456 7501
rect 8392 7452 8456 7467
rect 10050 7501 10114 7516
rect 10050 7467 10065 7501
rect 10099 7467 10114 7501
rect 10050 7452 10114 7467
rect -674 6394 -610 6409
rect -674 6360 -659 6394
rect -625 6360 -610 6394
rect -674 6345 -610 6360
rect 102 5091 166 5106
rect 102 5057 117 5091
rect 151 5057 166 5091
rect 102 5042 166 5057
rect 1760 5091 1824 5106
rect 1760 5057 1775 5091
rect 1809 5057 1824 5091
rect 1760 5042 1824 5057
rect 5076 5091 5140 5106
rect 5076 5057 5091 5091
rect 5125 5057 5140 5091
rect 5076 5042 5140 5057
rect 8392 5091 8456 5106
rect 8392 5057 8407 5091
rect 8441 5057 8456 5091
rect 8392 5042 8456 5057
rect 10050 5091 10114 5106
rect 10050 5057 10065 5091
rect 10099 5057 10114 5091
rect 10050 5042 10114 5057
rect -1831 4680 -1767 4695
rect -1831 4646 -1816 4680
rect -1782 4646 -1767 4680
rect -1831 4631 -1767 4646
rect 102 4168 166 4183
rect 102 4134 117 4168
rect 151 4134 166 4168
rect 102 4119 166 4134
rect 1760 4168 1824 4183
rect 1760 4134 1775 4168
rect 1809 4134 1824 4168
rect 1760 4119 1824 4134
rect 5076 4168 5140 4183
rect 5076 4134 5091 4168
rect 5125 4134 5140 4168
rect 5076 4119 5140 4134
rect 8392 4168 8456 4183
rect 8392 4134 8407 4168
rect 8441 4134 8456 4168
rect 8392 4119 8456 4134
rect 10050 4168 10114 4183
rect 10050 4134 10065 4168
rect 10099 4134 10114 4168
rect 10050 4119 10114 4134
rect -1831 3800 -1767 3815
rect -1831 3766 -1816 3800
rect -1782 3766 -1767 3800
rect -1831 3751 -1767 3766
rect 102 3288 166 3303
rect 102 3254 117 3288
rect 151 3254 166 3288
rect 102 3239 166 3254
rect 1760 3288 1824 3303
rect 1760 3254 1775 3288
rect 1809 3254 1824 3288
rect 1760 3239 1824 3254
rect 5076 3288 5140 3303
rect 5076 3254 5091 3288
rect 5125 3254 5140 3288
rect 5076 3239 5140 3254
rect 8392 3288 8456 3303
rect 8392 3254 8407 3288
rect 8441 3254 8456 3288
rect 8392 3239 8456 3254
rect 10050 3288 10114 3303
rect 10050 3254 10065 3288
rect 10099 3254 10114 3288
rect 10050 3239 10114 3254
rect 3418 2105 3482 2120
rect 3418 2071 3433 2105
rect 3467 2071 3482 2105
rect 3418 2056 3482 2071
rect 6734 2105 6798 2120
rect 6734 2071 6749 2105
rect 6783 2071 6798 2105
rect 6734 2056 6798 2071
rect 3418 17 3482 32
rect 3418 -17 3433 17
rect 3467 -17 3482 17
rect 3418 -32 3482 -17
rect 6734 16 6798 31
rect 6734 -18 6749 16
rect 6783 -18 6798 16
rect 6734 -33 6798 -18
<< viali >>
rect 117 7467 151 7501
rect 1775 7467 1809 7501
rect 5091 7467 5125 7501
rect 8407 7467 8441 7501
rect 10065 7467 10099 7501
rect -659 6360 -625 6394
rect 117 5057 151 5091
rect 1775 5057 1809 5091
rect 5091 5057 5125 5091
rect 8407 5057 8441 5091
rect 10065 5057 10099 5091
rect -1816 4646 -1782 4680
rect 117 4134 151 4168
rect 1775 4134 1809 4168
rect 5091 4134 5125 4168
rect 8407 4134 8441 4168
rect 10065 4134 10099 4168
rect -1816 3766 -1782 3800
rect 117 3254 151 3288
rect 1775 3254 1809 3288
rect 5091 3254 5125 3288
rect 8407 3254 8441 3288
rect 10065 3254 10099 3288
rect 3433 2071 3467 2105
rect 6749 2071 6783 2105
rect 3433 -17 3467 17
rect 6749 -18 6783 16
<< metal1 >>
rect 102 7510 166 7516
rect 102 7458 108 7510
rect 160 7458 166 7510
rect 102 7452 166 7458
rect 1760 7510 1824 7516
rect 1760 7458 1766 7510
rect 1818 7458 1824 7510
rect 1760 7452 1824 7458
rect 5076 7510 5140 7516
rect 5076 7458 5082 7510
rect 5134 7458 5140 7510
rect 5076 7452 5140 7458
rect 8392 7510 8456 7516
rect 8392 7458 8398 7510
rect 8450 7458 8456 7510
rect 8392 7452 8456 7458
rect 10050 7510 10114 7516
rect 10050 7458 10056 7510
rect 10108 7458 10114 7510
rect 10050 7452 10114 7458
rect 102 7336 166 7342
rect 102 7284 108 7336
rect 160 7284 166 7336
rect 102 7278 166 7284
rect 1760 7336 1824 7342
rect 1760 7284 1766 7336
rect 1818 7284 1824 7336
rect 1760 7278 1824 7284
rect 3418 7336 3482 7342
rect 3418 7284 3424 7336
rect 3476 7284 3482 7336
rect 3418 7278 3482 7284
rect 5076 7336 5140 7342
rect 5076 7284 5082 7336
rect 5134 7284 5140 7336
rect 5076 7278 5140 7284
rect 6734 7336 6798 7342
rect 6734 7284 6740 7336
rect 6792 7284 6798 7336
rect 6734 7278 6798 7284
rect 8392 7336 8456 7342
rect 8392 7284 8398 7336
rect 8450 7284 8456 7336
rect 8392 7278 8456 7284
rect 10050 7336 10114 7342
rect 10050 7284 10056 7336
rect 10108 7284 10114 7336
rect 10050 7278 10114 7284
rect 111 7227 157 7268
rect 3427 7227 3473 7268
rect 6743 7227 6789 7268
rect 10059 7227 10105 7268
rect 111 7181 167 7227
rect 3417 7181 3483 7227
rect 6733 7181 6799 7227
rect 10049 7181 10105 7227
rect 3427 7093 3473 7181
rect 6743 7093 6789 7181
rect 102 7087 166 7093
rect 102 7035 108 7087
rect 160 7035 166 7087
rect 102 7029 166 7035
rect 1760 7087 1824 7093
rect 1760 7035 1766 7087
rect 1818 7035 1824 7087
rect 1760 7029 1824 7035
rect 3418 7087 3482 7093
rect 3418 7035 3424 7087
rect 3476 7035 3482 7087
rect 3418 7029 3482 7035
rect 5076 7087 5140 7093
rect 5076 7035 5082 7087
rect 5134 7035 5140 7087
rect 5076 7029 5140 7035
rect 6734 7087 6798 7093
rect 6734 7035 6740 7087
rect 6792 7035 6798 7087
rect 6734 7029 6798 7035
rect 8392 7087 8456 7093
rect 8392 7035 8398 7087
rect 8450 7035 8456 7087
rect 8392 7029 8456 7035
rect 10050 7087 10114 7093
rect 10050 7035 10056 7087
rect 10108 7035 10114 7087
rect 10050 7029 10114 7035
rect 111 6978 157 7019
rect 3427 6978 3473 7029
rect 6743 6978 6789 7029
rect 10059 6978 10105 7019
rect 111 6932 167 6978
rect 3417 6932 3483 6978
rect 6733 6932 6799 6978
rect 10049 6932 10105 6978
rect 3427 6844 3473 6932
rect 6743 6844 6789 6932
rect 102 6838 166 6844
rect 102 6786 108 6838
rect 160 6786 166 6838
rect 102 6780 166 6786
rect 1760 6838 1824 6844
rect 1760 6786 1766 6838
rect 1818 6786 1824 6838
rect 1760 6780 1824 6786
rect 3418 6838 3482 6844
rect 3418 6786 3424 6838
rect 3476 6786 3482 6838
rect 3418 6780 3482 6786
rect 5076 6838 5140 6844
rect 5076 6786 5082 6838
rect 5134 6786 5140 6838
rect 5076 6780 5140 6786
rect 6734 6838 6798 6844
rect 6734 6786 6740 6838
rect 6792 6786 6798 6838
rect 6734 6780 6798 6786
rect 8392 6838 8456 6844
rect 8392 6786 8398 6838
rect 8450 6786 8456 6838
rect 8392 6780 8456 6786
rect 10050 6838 10114 6844
rect 10050 6786 10056 6838
rect 10108 6786 10114 6838
rect 10050 6780 10114 6786
rect 111 6729 157 6770
rect 3427 6729 3473 6780
rect 6743 6729 6789 6780
rect 10059 6729 10105 6770
rect 111 6683 167 6729
rect 3417 6683 3483 6729
rect 6733 6683 6799 6729
rect 10049 6683 10105 6729
rect 3427 6595 3473 6683
rect 6743 6595 6789 6683
rect 102 6589 166 6595
rect 102 6537 108 6589
rect 160 6537 166 6589
rect 102 6531 166 6537
rect 1760 6589 1824 6595
rect 1760 6537 1766 6589
rect 1818 6537 1824 6589
rect 1760 6531 1824 6537
rect 3418 6589 3482 6595
rect 3418 6537 3424 6589
rect 3476 6537 3482 6589
rect 3418 6531 3482 6537
rect 5076 6589 5140 6595
rect 5076 6537 5082 6589
rect 5134 6537 5140 6589
rect 5076 6531 5140 6537
rect 6734 6589 6798 6595
rect 6734 6537 6740 6589
rect 6792 6537 6798 6589
rect 6734 6531 6798 6537
rect 8392 6589 8456 6595
rect 8392 6537 8398 6589
rect 8450 6537 8456 6589
rect 8392 6531 8456 6537
rect 10050 6589 10114 6595
rect 10050 6537 10056 6589
rect 10108 6537 10114 6589
rect 10050 6531 10114 6537
rect 111 6480 157 6521
rect 3427 6480 3473 6531
rect 6743 6480 6789 6531
rect 10059 6480 10105 6521
rect 111 6434 167 6480
rect 3417 6434 3483 6480
rect 6733 6434 6799 6480
rect 10049 6434 10105 6480
rect -1035 6416 -971 6422
rect -1035 6364 -1029 6416
rect -977 6364 -971 6416
rect -1035 6358 -971 6364
rect -674 6403 -610 6409
rect -674 6351 -668 6403
rect -616 6351 -610 6403
rect -674 6345 -610 6351
rect 102 6340 166 6346
rect 102 6288 108 6340
rect 160 6288 166 6340
rect 102 6282 166 6288
rect 1760 6340 1824 6346
rect 1760 6288 1766 6340
rect 1818 6288 1824 6340
rect 1760 6282 1824 6288
rect 3418 6340 3482 6346
rect 3418 6288 3424 6340
rect 3476 6288 3482 6340
rect 3418 6282 3482 6288
rect 5076 6340 5140 6346
rect 5076 6288 5082 6340
rect 5134 6288 5140 6340
rect 5076 6282 5140 6288
rect 6734 6340 6798 6346
rect 6734 6288 6740 6340
rect 6792 6288 6798 6340
rect 6734 6282 6798 6288
rect 8392 6340 8456 6346
rect 8392 6288 8398 6340
rect 8450 6288 8456 6340
rect 8392 6282 8456 6288
rect 10050 6340 10114 6346
rect 10050 6288 10056 6340
rect 10108 6288 10114 6340
rect 10050 6282 10114 6288
rect 111 6231 157 6272
rect 4300 6234 4364 6240
rect 111 6185 167 6231
rect 3417 6185 3483 6231
rect 4300 6182 4306 6234
rect 4358 6182 4364 6234
rect 4300 6176 4364 6182
rect 5956 6234 6020 6240
rect 5956 6182 5962 6234
rect 6014 6182 6020 6234
rect 10059 6231 10105 6272
rect 6733 6185 6799 6231
rect 10049 6185 10105 6231
rect 5956 6176 6020 6182
rect 102 6091 166 6097
rect 102 6039 108 6091
rect 160 6039 166 6091
rect 102 6033 166 6039
rect 1760 6091 1824 6097
rect 1760 6039 1766 6091
rect 1818 6039 1824 6091
rect 1760 6033 1824 6039
rect 3418 6091 3482 6097
rect 3418 6039 3424 6091
rect 3476 6039 3482 6091
rect 3418 6033 3482 6039
rect 5076 6091 5140 6097
rect 5076 6039 5082 6091
rect 5134 6039 5140 6091
rect 5076 6033 5140 6039
rect 6734 6091 6798 6097
rect 6734 6039 6740 6091
rect 6792 6039 6798 6091
rect 6734 6033 6798 6039
rect 8392 6091 8456 6097
rect 8392 6039 8398 6091
rect 8450 6039 8456 6091
rect 8392 6033 8456 6039
rect 10050 6091 10114 6097
rect 10050 6039 10056 6091
rect 10108 6039 10114 6091
rect 10050 6033 10114 6039
rect 111 5982 157 6023
rect 4300 5985 4364 5991
rect 111 5936 167 5982
rect 3417 5936 3483 5982
rect 4300 5933 4306 5985
rect 4358 5933 4364 5985
rect 4300 5927 4364 5933
rect 5956 5985 6020 5991
rect 5956 5933 5962 5985
rect 6014 5933 6020 5985
rect 10059 5982 10105 6023
rect 6733 5936 6799 5982
rect 10049 5936 10105 5982
rect 5956 5927 6020 5933
rect 102 5842 166 5848
rect 102 5790 108 5842
rect 160 5790 166 5842
rect 102 5784 166 5790
rect 1760 5842 1824 5848
rect 1760 5790 1766 5842
rect 1818 5790 1824 5842
rect 1760 5784 1824 5790
rect 3418 5842 3482 5848
rect 3418 5790 3424 5842
rect 3476 5790 3482 5842
rect 3418 5784 3482 5790
rect 5076 5842 5140 5848
rect 5076 5790 5082 5842
rect 5134 5790 5140 5842
rect 5076 5784 5140 5790
rect 6734 5842 6798 5848
rect 6734 5790 6740 5842
rect 6792 5790 6798 5842
rect 6734 5784 6798 5790
rect 8392 5842 8456 5848
rect 8392 5790 8398 5842
rect 8450 5790 8456 5842
rect 8392 5784 8456 5790
rect 10050 5842 10114 5848
rect 10050 5790 10056 5842
rect 10108 5790 10114 5842
rect 10050 5784 10114 5790
rect 111 5733 157 5774
rect 4300 5736 4364 5742
rect 111 5687 167 5733
rect 3417 5687 3483 5733
rect 4300 5684 4306 5736
rect 4358 5684 4364 5736
rect 4300 5678 4364 5684
rect 5956 5736 6020 5742
rect 5956 5684 5962 5736
rect 6014 5684 6020 5736
rect 10059 5733 10105 5774
rect 6733 5687 6799 5733
rect 10049 5687 10105 5733
rect 5956 5678 6020 5684
rect 102 5593 166 5599
rect 102 5541 108 5593
rect 160 5541 166 5593
rect 102 5535 166 5541
rect 1760 5593 1824 5599
rect 1760 5541 1766 5593
rect 1818 5541 1824 5593
rect 1760 5535 1824 5541
rect 3418 5593 3482 5599
rect 3418 5541 3424 5593
rect 3476 5541 3482 5593
rect 3418 5535 3482 5541
rect 5076 5593 5140 5599
rect 5076 5541 5082 5593
rect 5134 5541 5140 5593
rect 5076 5535 5140 5541
rect 6734 5593 6798 5599
rect 6734 5541 6740 5593
rect 6792 5541 6798 5593
rect 6734 5535 6798 5541
rect 8392 5593 8456 5599
rect 8392 5541 8398 5593
rect 8450 5541 8456 5593
rect 8392 5535 8456 5541
rect 10050 5593 10114 5599
rect 10050 5541 10056 5593
rect 10108 5541 10114 5593
rect 10050 5535 10114 5541
rect 111 5484 157 5525
rect 4300 5487 4364 5493
rect 111 5438 167 5484
rect 3417 5438 3483 5484
rect 4300 5435 4306 5487
rect 4358 5435 4364 5487
rect 4300 5429 4364 5435
rect 5956 5487 6020 5493
rect 5956 5435 5962 5487
rect 6014 5435 6020 5487
rect 10059 5484 10105 5525
rect 6733 5438 6799 5484
rect 10049 5438 10105 5484
rect 5956 5429 6020 5435
rect 102 5344 166 5350
rect 102 5292 108 5344
rect 160 5292 166 5344
rect 102 5286 166 5292
rect 1760 5344 1824 5350
rect 1760 5292 1766 5344
rect 1818 5292 1824 5344
rect 1760 5286 1824 5292
rect 3418 5344 3482 5350
rect 3418 5292 3424 5344
rect 3476 5292 3482 5344
rect 3418 5286 3482 5292
rect 5076 5344 5140 5350
rect 5076 5292 5082 5344
rect 5134 5292 5140 5344
rect 5076 5286 5140 5292
rect 6734 5344 6798 5350
rect 6734 5292 6740 5344
rect 6792 5292 6798 5344
rect 6734 5286 6798 5292
rect 8392 5344 8456 5350
rect 8392 5292 8398 5344
rect 8450 5292 8456 5344
rect 8392 5286 8456 5292
rect 10050 5344 10114 5350
rect 10050 5292 10056 5344
rect 10108 5292 10114 5344
rect 10050 5286 10114 5292
rect 111 5235 157 5276
rect 4300 5238 4364 5244
rect 111 5189 167 5235
rect 3417 5189 3483 5235
rect 4300 5186 4306 5238
rect 4358 5186 4364 5238
rect 4300 5180 4364 5186
rect 5956 5238 6020 5244
rect 5956 5186 5962 5238
rect 6014 5186 6020 5238
rect 10059 5235 10105 5276
rect 6733 5189 6799 5235
rect 10049 5189 10105 5235
rect 5956 5180 6020 5186
rect 102 5100 166 5106
rect 102 5048 108 5100
rect 160 5048 166 5100
rect 102 5042 166 5048
rect 1760 5100 1824 5106
rect 1760 5048 1766 5100
rect 1818 5048 1824 5100
rect 1760 5042 1824 5048
rect 5076 5100 5140 5106
rect 5076 5048 5082 5100
rect 5134 5048 5140 5100
rect 5076 5042 5140 5048
rect 8392 5100 8456 5106
rect 8392 5048 8398 5100
rect 8450 5048 8456 5100
rect 8392 5042 8456 5048
rect 10050 5100 10114 5106
rect 10050 5048 10056 5100
rect 10108 5048 10114 5100
rect 10050 5042 10114 5048
rect 102 4937 166 4943
rect 102 4885 108 4937
rect 160 4885 166 4937
rect 102 4879 166 4885
rect 1760 4937 1824 4943
rect 1760 4885 1766 4937
rect 1818 4885 1824 4937
rect 1760 4879 1824 4885
rect 5076 4937 5140 4943
rect 5076 4885 5082 4937
rect 5134 4885 5140 4937
rect 5076 4879 5140 4885
rect 8392 4937 8456 4943
rect 8392 4885 8398 4937
rect 8450 4885 8456 4937
rect 8392 4879 8456 4885
rect 10050 4937 10114 4943
rect 10050 4885 10056 4937
rect 10108 4885 10114 4937
rect 10050 4879 10114 4885
rect 3418 4807 3482 4813
rect 3418 4755 3424 4807
rect 3476 4755 3482 4807
rect 3418 4749 3482 4755
rect 6734 4807 6798 4813
rect 6734 4755 6740 4807
rect 6792 4755 6798 4807
rect 6734 4749 6798 4755
rect 111 4702 157 4743
rect 4300 4705 4364 4711
rect -1831 4689 -1767 4695
rect -1831 4637 -1825 4689
rect -1773 4637 -1767 4689
rect 111 4656 167 4702
rect 3417 4656 3483 4702
rect 4300 4653 4306 4705
rect 4358 4653 4364 4705
rect 4300 4647 4364 4653
rect 5956 4705 6020 4711
rect 5956 4653 5962 4705
rect 6014 4653 6020 4705
rect 10059 4702 10105 4743
rect 6733 4656 6799 4702
rect 10049 4656 10105 4702
rect 5956 4647 6020 4653
rect -1831 4631 -1767 4637
rect -1831 4458 -1767 4464
rect -1831 4406 -1825 4458
rect -1773 4406 -1767 4458
rect -1831 4400 -1767 4406
rect 102 4177 166 4183
rect 102 4125 108 4177
rect 160 4125 166 4177
rect 102 4119 166 4125
rect 1760 4177 1824 4183
rect 1760 4125 1766 4177
rect 1818 4125 1824 4177
rect 1760 4119 1824 4125
rect 5076 4177 5140 4183
rect 5076 4125 5082 4177
rect 5134 4125 5140 4177
rect 5076 4119 5140 4125
rect 8392 4177 8456 4183
rect 8392 4125 8398 4177
rect 8450 4125 8456 4177
rect 8392 4119 8456 4125
rect 10050 4177 10114 4183
rect 10050 4125 10056 4177
rect 10108 4125 10114 4177
rect 10050 4119 10114 4125
rect -1831 4102 -1767 4108
rect -1831 4050 -1825 4102
rect -1773 4050 -1767 4102
rect -1831 4044 -1767 4050
rect 108 3990 167 4036
rect 3417 3990 3483 4036
rect 5075 3990 5141 4036
rect 6733 3990 6799 4036
rect 10049 3990 10108 4036
rect 108 3952 160 3990
rect 3427 3952 3473 3990
rect 10056 3952 10108 3990
rect 102 3946 166 3952
rect 102 3894 108 3946
rect 160 3894 166 3946
rect 102 3888 166 3894
rect 1760 3946 1824 3952
rect 1760 3894 1766 3946
rect 1818 3894 1824 3946
rect 1760 3888 1824 3894
rect 3418 3946 3482 3952
rect 3418 3894 3424 3946
rect 3476 3894 3482 3946
rect 3418 3888 3482 3894
rect 5076 3946 5140 3952
rect 5076 3894 5082 3946
rect 5134 3894 5140 3946
rect 5076 3888 5140 3894
rect 6734 3946 6798 3952
rect 6734 3894 6740 3946
rect 6792 3894 6798 3946
rect 6734 3888 6798 3894
rect 8392 3946 8456 3952
rect 8392 3894 8398 3946
rect 8450 3894 8456 3946
rect 8392 3888 8456 3894
rect 10050 3946 10114 3952
rect 10050 3894 10056 3946
rect 10108 3894 10114 3946
rect 10050 3888 10114 3894
rect -1831 3809 -1767 3815
rect -1831 3757 -1825 3809
rect -1773 3757 -1767 3809
rect -1831 3751 -1767 3757
rect 108 3634 167 3680
rect 3417 3634 3483 3680
rect 5075 3634 5141 3680
rect 6733 3634 6799 3680
rect 10049 3634 10108 3680
rect 108 3596 160 3634
rect 3427 3596 3473 3634
rect 10056 3596 10108 3634
rect 102 3590 166 3596
rect 102 3538 108 3590
rect 160 3538 166 3590
rect 102 3532 166 3538
rect 1760 3590 1824 3596
rect 1760 3538 1766 3590
rect 1818 3538 1824 3590
rect 1760 3532 1824 3538
rect 3418 3590 3482 3596
rect 3418 3538 3424 3590
rect 3476 3538 3482 3590
rect 3418 3532 3482 3538
rect 5076 3590 5140 3596
rect 5076 3538 5082 3590
rect 5134 3538 5140 3590
rect 5076 3532 5140 3538
rect 8392 3590 8456 3596
rect 8392 3538 8398 3590
rect 8450 3538 8456 3590
rect 8392 3532 8456 3538
rect 10050 3590 10114 3596
rect 10050 3538 10056 3590
rect 10108 3538 10114 3590
rect 10050 3532 10114 3538
rect 6734 3466 6798 3472
rect 6734 3414 6740 3466
rect 6792 3414 6798 3466
rect 6734 3408 6798 3414
rect 102 3297 166 3303
rect 102 3245 108 3297
rect 160 3245 166 3297
rect 102 3239 166 3245
rect 1760 3297 1824 3303
rect 1760 3245 1766 3297
rect 1818 3245 1824 3297
rect 1760 3239 1824 3245
rect 5076 3297 5140 3303
rect 5076 3245 5082 3297
rect 5134 3245 5140 3297
rect 5076 3239 5140 3245
rect 8392 3297 8456 3303
rect 8392 3245 8398 3297
rect 8450 3245 8456 3297
rect 8392 3239 8456 3245
rect 10050 3297 10114 3303
rect 10050 3245 10056 3297
rect 10108 3245 10114 3297
rect 10050 3239 10114 3245
rect 3418 2114 3482 2120
rect 3418 2062 3424 2114
rect 3476 2062 3482 2114
rect 3418 2056 3482 2062
rect 6734 2114 6798 2120
rect 6734 2062 6740 2114
rect 6792 2062 6798 2114
rect 6734 2056 6798 2062
rect 3138 1976 3202 1982
rect 3138 1924 3144 1976
rect 3196 1924 3202 1976
rect 3138 1918 3202 1924
rect 4725 1976 4789 1982
rect 4725 1924 4731 1976
rect 4783 1924 4789 1976
rect 6957 1976 7021 1982
rect 5075 1927 5141 1973
rect 4725 1918 4789 1924
rect 6957 1924 6963 1976
rect 7015 1924 7021 1976
rect 6957 1918 7021 1924
rect 102 1827 108 1879
rect 160 1827 166 1879
rect 1760 1827 1766 1879
rect 1818 1827 1824 1879
rect 3418 1827 3424 1879
rect 3476 1827 3482 1879
rect 5076 1827 5082 1879
rect 5134 1827 5140 1879
rect 6734 1827 6740 1879
rect 6792 1827 6798 1879
rect 8392 1827 8398 1879
rect 8450 1827 8456 1879
rect 10050 1827 10056 1879
rect 10108 1827 10114 1879
rect 3138 1736 3202 1742
rect 3138 1684 3144 1736
rect 3196 1684 3202 1736
rect 3138 1678 3202 1684
rect 4725 1736 4789 1742
rect 4725 1684 4731 1736
rect 4783 1684 4789 1736
rect 6957 1736 7021 1742
rect 5075 1687 5141 1733
rect 4725 1678 4789 1684
rect 6957 1684 6963 1736
rect 7015 1684 7021 1736
rect 6957 1678 7021 1684
rect 102 1587 108 1639
rect 160 1587 166 1639
rect 1760 1587 1766 1639
rect 1818 1587 1824 1639
rect 3418 1587 3424 1639
rect 3476 1587 3482 1639
rect 5076 1587 5082 1639
rect 5134 1587 5140 1639
rect 6734 1587 6740 1639
rect 6792 1587 6798 1639
rect 8392 1587 8398 1639
rect 8450 1587 8456 1639
rect 10050 1587 10056 1639
rect 10108 1587 10114 1639
rect 3138 1496 3202 1502
rect 3138 1444 3144 1496
rect 3196 1444 3202 1496
rect 3138 1438 3202 1444
rect 4725 1496 4789 1502
rect 4725 1444 4731 1496
rect 4783 1444 4789 1496
rect 6957 1496 7021 1502
rect 5075 1447 5141 1493
rect 4725 1438 4789 1444
rect 6957 1444 6963 1496
rect 7015 1444 7021 1496
rect 6957 1438 7021 1444
rect 102 1347 108 1399
rect 160 1347 166 1399
rect 1760 1347 1766 1399
rect 1818 1347 1824 1399
rect 3418 1347 3424 1399
rect 3476 1347 3482 1399
rect 5076 1347 5082 1399
rect 5134 1347 5140 1399
rect 6734 1347 6740 1399
rect 6792 1347 6798 1399
rect 8392 1347 8398 1399
rect 8450 1347 8456 1399
rect 10050 1347 10056 1399
rect 10108 1347 10114 1399
rect 3138 1256 3202 1262
rect 3138 1204 3144 1256
rect 3196 1204 3202 1256
rect 3138 1198 3202 1204
rect 4725 1256 4789 1262
rect 4725 1204 4731 1256
rect 4783 1204 4789 1256
rect 6957 1256 7021 1262
rect 5075 1207 5141 1253
rect 4725 1198 4789 1204
rect 6957 1204 6963 1256
rect 7015 1204 7021 1256
rect 6957 1198 7021 1204
rect 102 1107 108 1159
rect 160 1107 166 1159
rect 1760 1107 1766 1159
rect 1818 1107 1824 1159
rect 3418 1107 3424 1159
rect 3476 1107 3482 1159
rect 5076 1107 5082 1159
rect 5134 1107 5140 1159
rect 6734 1107 6740 1159
rect 6792 1107 6798 1159
rect 8392 1107 8398 1159
rect 8450 1107 8456 1159
rect 10050 1107 10056 1159
rect 10108 1107 10114 1159
rect 3138 1016 3202 1022
rect 3138 964 3144 1016
rect 3196 964 3202 1016
rect 3138 958 3202 964
rect 4725 1016 4789 1022
rect 4725 964 4731 1016
rect 4783 964 4789 1016
rect 6957 1016 7021 1022
rect 5075 967 5141 1013
rect 4725 958 4789 964
rect 6957 964 6963 1016
rect 7015 964 7021 1016
rect 6957 958 7021 964
rect 102 867 108 919
rect 160 867 166 919
rect 1760 867 1766 919
rect 1818 867 1824 919
rect 3418 867 3424 919
rect 3476 867 3482 919
rect 5076 867 5082 919
rect 5134 867 5140 919
rect 6734 867 6740 919
rect 6792 867 6798 919
rect 8392 867 8398 919
rect 8450 867 8456 919
rect 10050 867 10056 919
rect 10108 867 10114 919
rect 3138 776 3202 782
rect 3138 724 3144 776
rect 3196 724 3202 776
rect 3138 718 3202 724
rect 4725 776 4789 782
rect 4725 724 4731 776
rect 4783 724 4789 776
rect 6957 776 7021 782
rect 5075 727 5141 773
rect 4725 718 4789 724
rect 6957 724 6963 776
rect 7015 724 7021 776
rect 6957 718 7021 724
rect 102 627 108 679
rect 160 627 166 679
rect 1760 627 1766 679
rect 1818 627 1824 679
rect 3418 627 3424 679
rect 3476 627 3482 679
rect 5076 627 5082 679
rect 5134 627 5140 679
rect 6734 627 6740 679
rect 6792 627 6798 679
rect 8392 627 8398 679
rect 8450 627 8456 679
rect 10050 627 10056 679
rect 10108 627 10114 679
rect 3138 536 3202 542
rect 3138 484 3144 536
rect 3196 484 3202 536
rect 3138 478 3202 484
rect 4725 536 4789 542
rect 4725 484 4731 536
rect 4783 484 4789 536
rect 6957 536 7021 542
rect 5075 487 5141 533
rect 4725 478 4789 484
rect 6957 484 6963 536
rect 7015 484 7021 536
rect 6957 478 7021 484
rect 102 387 108 439
rect 160 387 166 439
rect 1760 387 1766 439
rect 1818 387 1824 439
rect 3418 387 3424 439
rect 3476 387 3482 439
rect 5076 387 5082 439
rect 5134 387 5140 439
rect 6734 387 6740 439
rect 6792 387 6798 439
rect 8392 387 8398 439
rect 8450 387 8456 439
rect 10050 387 10056 439
rect 10108 387 10114 439
rect 3138 296 3202 302
rect 3138 244 3144 296
rect 3196 244 3202 296
rect 3138 238 3202 244
rect 4725 296 4789 302
rect 4725 244 4731 296
rect 4783 244 4789 296
rect 6957 296 7021 302
rect 5075 247 5141 293
rect 4725 238 4789 244
rect 6957 244 6963 296
rect 7015 244 7021 296
rect 6957 238 7021 244
rect 102 147 108 199
rect 160 147 166 199
rect 1760 147 1766 199
rect 1818 147 1824 199
rect 3418 147 3424 199
rect 3476 147 3482 199
rect 5076 147 5082 199
rect 5134 147 5140 199
rect 6734 147 6740 199
rect 6792 147 6798 199
rect 8392 147 8398 199
rect 8450 147 8456 199
rect 10050 147 10056 199
rect 10108 147 10114 199
rect 3418 26 3482 32
rect 3418 -26 3424 26
rect 3476 -26 3482 26
rect 3418 -32 3482 -26
rect 6734 25 6798 31
rect 6734 -27 6740 25
rect 6792 -27 6798 25
rect 6734 -33 6798 -27
<< via1 >>
rect 108 7501 160 7510
rect 108 7467 117 7501
rect 117 7467 151 7501
rect 151 7467 160 7501
rect 108 7458 160 7467
rect 1766 7501 1818 7510
rect 1766 7467 1775 7501
rect 1775 7467 1809 7501
rect 1809 7467 1818 7501
rect 1766 7458 1818 7467
rect 5082 7501 5134 7510
rect 5082 7467 5091 7501
rect 5091 7467 5125 7501
rect 5125 7467 5134 7501
rect 5082 7458 5134 7467
rect 8398 7501 8450 7510
rect 8398 7467 8407 7501
rect 8407 7467 8441 7501
rect 8441 7467 8450 7501
rect 8398 7458 8450 7467
rect 10056 7501 10108 7510
rect 10056 7467 10065 7501
rect 10065 7467 10099 7501
rect 10099 7467 10108 7501
rect 10056 7458 10108 7467
rect 108 7284 160 7336
rect 1766 7284 1818 7336
rect 3424 7284 3476 7336
rect 5082 7284 5134 7336
rect 6740 7284 6792 7336
rect 8398 7284 8450 7336
rect 10056 7284 10108 7336
rect 108 7035 160 7087
rect 1766 7035 1818 7087
rect 3424 7035 3476 7087
rect 5082 7035 5134 7087
rect 6740 7035 6792 7087
rect 8398 7035 8450 7087
rect 10056 7035 10108 7087
rect 108 6786 160 6838
rect 1766 6786 1818 6838
rect 3424 6786 3476 6838
rect 5082 6786 5134 6838
rect 6740 6786 6792 6838
rect 8398 6786 8450 6838
rect 10056 6786 10108 6838
rect 108 6537 160 6589
rect 1766 6537 1818 6589
rect 3424 6537 3476 6589
rect 5082 6537 5134 6589
rect 6740 6537 6792 6589
rect 8398 6537 8450 6589
rect 10056 6537 10108 6589
rect -1029 6364 -977 6416
rect -668 6394 -616 6403
rect -668 6360 -659 6394
rect -659 6360 -625 6394
rect -625 6360 -616 6394
rect -668 6351 -616 6360
rect 108 6288 160 6340
rect 1766 6288 1818 6340
rect 3424 6288 3476 6340
rect 5082 6288 5134 6340
rect 6740 6288 6792 6340
rect 8398 6288 8450 6340
rect 10056 6288 10108 6340
rect 4306 6182 4358 6234
rect 5962 6182 6014 6234
rect 108 6039 160 6091
rect 1766 6039 1818 6091
rect 3424 6039 3476 6091
rect 5082 6039 5134 6091
rect 6740 6039 6792 6091
rect 8398 6039 8450 6091
rect 10056 6039 10108 6091
rect 4306 5933 4358 5985
rect 5962 5933 6014 5985
rect 108 5790 160 5842
rect 1766 5790 1818 5842
rect 3424 5790 3476 5842
rect 5082 5790 5134 5842
rect 6740 5790 6792 5842
rect 8398 5790 8450 5842
rect 10056 5790 10108 5842
rect 4306 5684 4358 5736
rect 5962 5684 6014 5736
rect 108 5541 160 5593
rect 1766 5541 1818 5593
rect 3424 5541 3476 5593
rect 5082 5541 5134 5593
rect 6740 5541 6792 5593
rect 8398 5541 8450 5593
rect 10056 5541 10108 5593
rect 4306 5435 4358 5487
rect 5962 5435 6014 5487
rect 108 5292 160 5344
rect 1766 5292 1818 5344
rect 3424 5292 3476 5344
rect 5082 5292 5134 5344
rect 6740 5292 6792 5344
rect 8398 5292 8450 5344
rect 10056 5292 10108 5344
rect 4306 5186 4358 5238
rect 5962 5186 6014 5238
rect 108 5091 160 5100
rect 108 5057 117 5091
rect 117 5057 151 5091
rect 151 5057 160 5091
rect 108 5048 160 5057
rect 1766 5091 1818 5100
rect 1766 5057 1775 5091
rect 1775 5057 1809 5091
rect 1809 5057 1818 5091
rect 1766 5048 1818 5057
rect 5082 5091 5134 5100
rect 5082 5057 5091 5091
rect 5091 5057 5125 5091
rect 5125 5057 5134 5091
rect 5082 5048 5134 5057
rect 8398 5091 8450 5100
rect 8398 5057 8407 5091
rect 8407 5057 8441 5091
rect 8441 5057 8450 5091
rect 8398 5048 8450 5057
rect 10056 5091 10108 5100
rect 10056 5057 10065 5091
rect 10065 5057 10099 5091
rect 10099 5057 10108 5091
rect 10056 5048 10108 5057
rect 108 4885 160 4937
rect 1766 4885 1818 4937
rect 5082 4885 5134 4937
rect 8398 4885 8450 4937
rect 10056 4885 10108 4937
rect 3424 4755 3476 4807
rect 6740 4755 6792 4807
rect -1825 4680 -1773 4689
rect -1825 4646 -1816 4680
rect -1816 4646 -1782 4680
rect -1782 4646 -1773 4680
rect -1825 4637 -1773 4646
rect 4306 4653 4358 4705
rect 5962 4653 6014 4705
rect -1825 4406 -1773 4458
rect 108 4168 160 4177
rect 108 4134 117 4168
rect 117 4134 151 4168
rect 151 4134 160 4168
rect 108 4125 160 4134
rect 1766 4168 1818 4177
rect 1766 4134 1775 4168
rect 1775 4134 1809 4168
rect 1809 4134 1818 4168
rect 1766 4125 1818 4134
rect 5082 4168 5134 4177
rect 5082 4134 5091 4168
rect 5091 4134 5125 4168
rect 5125 4134 5134 4168
rect 5082 4125 5134 4134
rect 8398 4168 8450 4177
rect 8398 4134 8407 4168
rect 8407 4134 8441 4168
rect 8441 4134 8450 4168
rect 8398 4125 8450 4134
rect 10056 4168 10108 4177
rect 10056 4134 10065 4168
rect 10065 4134 10099 4168
rect 10099 4134 10108 4168
rect 10056 4125 10108 4134
rect -1825 4050 -1773 4102
rect 108 3894 160 3946
rect 1766 3894 1818 3946
rect 3424 3894 3476 3946
rect 5082 3894 5134 3946
rect 6740 3894 6792 3946
rect 8398 3894 8450 3946
rect 10056 3894 10108 3946
rect -1825 3800 -1773 3809
rect -1825 3766 -1816 3800
rect -1816 3766 -1782 3800
rect -1782 3766 -1773 3800
rect -1825 3757 -1773 3766
rect 108 3538 160 3590
rect 1766 3538 1818 3590
rect 3424 3538 3476 3590
rect 5082 3538 5134 3590
rect 8398 3538 8450 3590
rect 10056 3538 10108 3590
rect 6740 3414 6792 3466
rect 108 3288 160 3297
rect 108 3254 117 3288
rect 117 3254 151 3288
rect 151 3254 160 3288
rect 108 3245 160 3254
rect 1766 3288 1818 3297
rect 1766 3254 1775 3288
rect 1775 3254 1809 3288
rect 1809 3254 1818 3288
rect 1766 3245 1818 3254
rect 5082 3288 5134 3297
rect 5082 3254 5091 3288
rect 5091 3254 5125 3288
rect 5125 3254 5134 3288
rect 5082 3245 5134 3254
rect 8398 3288 8450 3297
rect 8398 3254 8407 3288
rect 8407 3254 8441 3288
rect 8441 3254 8450 3288
rect 8398 3245 8450 3254
rect 10056 3288 10108 3297
rect 10056 3254 10065 3288
rect 10065 3254 10099 3288
rect 10099 3254 10108 3288
rect 10056 3245 10108 3254
rect 3424 2105 3476 2114
rect 3424 2071 3433 2105
rect 3433 2071 3467 2105
rect 3467 2071 3476 2105
rect 3424 2062 3476 2071
rect 6740 2105 6792 2114
rect 6740 2071 6749 2105
rect 6749 2071 6783 2105
rect 6783 2071 6792 2105
rect 6740 2062 6792 2071
rect 3144 1924 3196 1976
rect 4731 1924 4783 1976
rect 6963 1924 7015 1976
rect 108 1827 160 1879
rect 1766 1827 1818 1879
rect 3424 1827 3476 1879
rect 5082 1827 5134 1879
rect 6740 1827 6792 1879
rect 8398 1827 8450 1879
rect 10056 1827 10108 1879
rect 3144 1684 3196 1736
rect 4731 1684 4783 1736
rect 6963 1684 7015 1736
rect 108 1587 160 1639
rect 1766 1587 1818 1639
rect 3424 1587 3476 1639
rect 5082 1587 5134 1639
rect 6740 1587 6792 1639
rect 8398 1587 8450 1639
rect 10056 1587 10108 1639
rect 3144 1444 3196 1496
rect 4731 1444 4783 1496
rect 6963 1444 7015 1496
rect 108 1347 160 1399
rect 1766 1347 1818 1399
rect 3424 1347 3476 1399
rect 5082 1347 5134 1399
rect 6740 1347 6792 1399
rect 8398 1347 8450 1399
rect 10056 1347 10108 1399
rect 3144 1204 3196 1256
rect 4731 1204 4783 1256
rect 6963 1204 7015 1256
rect 108 1107 160 1159
rect 1766 1107 1818 1159
rect 3424 1107 3476 1159
rect 5082 1107 5134 1159
rect 6740 1107 6792 1159
rect 8398 1107 8450 1159
rect 10056 1107 10108 1159
rect 3144 964 3196 1016
rect 4731 964 4783 1016
rect 6963 964 7015 1016
rect 108 867 160 919
rect 1766 867 1818 919
rect 3424 867 3476 919
rect 5082 867 5134 919
rect 6740 867 6792 919
rect 8398 867 8450 919
rect 10056 867 10108 919
rect 3144 724 3196 776
rect 4731 724 4783 776
rect 6963 724 7015 776
rect 108 627 160 679
rect 1766 627 1818 679
rect 3424 627 3476 679
rect 5082 627 5134 679
rect 6740 627 6792 679
rect 8398 627 8450 679
rect 10056 627 10108 679
rect 3144 484 3196 536
rect 4731 484 4783 536
rect 6963 484 7015 536
rect 108 387 160 439
rect 1766 387 1818 439
rect 3424 387 3476 439
rect 5082 387 5134 439
rect 6740 387 6792 439
rect 8398 387 8450 439
rect 10056 387 10108 439
rect 3144 244 3196 296
rect 4731 244 4783 296
rect 6963 244 7015 296
rect 108 147 160 199
rect 1766 147 1818 199
rect 3424 147 3476 199
rect 5082 147 5134 199
rect 6740 147 6792 199
rect 8398 147 8450 199
rect 10056 147 10108 199
rect 3424 17 3476 26
rect 3424 -17 3433 17
rect 3433 -17 3467 17
rect 3467 -17 3476 17
rect 3424 -26 3476 -17
rect 6740 16 6792 25
rect 6740 -18 6749 16
rect 6749 -18 6783 16
rect 6783 -18 6792 16
rect 6740 -27 6792 -18
<< metal2 >>
rect 102 7510 166 7516
rect 102 7458 108 7510
rect 160 7458 166 7510
rect 102 7336 166 7458
rect 102 7284 108 7336
rect 160 7284 166 7336
rect 102 7087 166 7284
rect 102 7035 108 7087
rect 160 7035 166 7087
rect 102 6838 166 7035
rect 102 6786 108 6838
rect 160 6786 166 6838
rect 102 6589 166 6786
rect 102 6537 108 6589
rect 160 6537 166 6589
rect -1035 6416 -971 6422
rect -1035 6364 -1029 6416
rect -977 6364 -971 6416
rect -1035 6358 -971 6364
rect -674 6403 -610 6409
rect -674 6351 -668 6403
rect -616 6351 -610 6403
rect -674 6345 -610 6351
rect 102 6340 166 6537
rect 102 6288 108 6340
rect 160 6288 166 6340
rect -1039 6252 -965 6261
rect -1039 6196 -1030 6252
rect -974 6196 -965 6252
rect -1039 6187 -965 6196
rect 102 6091 166 6288
rect 102 6039 108 6091
rect 160 6039 166 6091
rect 102 5842 166 6039
rect 102 5790 108 5842
rect 160 5790 166 5842
rect 102 5593 166 5790
rect 102 5541 108 5593
rect 160 5541 166 5593
rect 102 5344 166 5541
rect 102 5292 108 5344
rect 160 5292 166 5344
rect 102 5100 166 5292
rect 102 5048 108 5100
rect 160 5048 166 5100
rect 102 4937 166 5048
rect 102 4885 108 4937
rect 160 4885 166 4937
rect 102 4879 166 4885
rect 1760 7510 1824 7516
rect 1760 7458 1766 7510
rect 1818 7458 1824 7510
rect 1760 7336 1824 7458
rect 5076 7510 5140 7516
rect 5076 7458 5082 7510
rect 5134 7458 5140 7510
rect 1760 7284 1766 7336
rect 1818 7284 1824 7336
rect 1760 7087 1824 7284
rect 1760 7035 1766 7087
rect 1818 7035 1824 7087
rect 1760 6838 1824 7035
rect 1760 6786 1766 6838
rect 1818 6786 1824 6838
rect 1760 6589 1824 6786
rect 1760 6537 1766 6589
rect 1818 6537 1824 6589
rect 1760 6340 1824 6537
rect 1760 6288 1766 6340
rect 1818 6288 1824 6340
rect 1760 6091 1824 6288
rect 1760 6039 1766 6091
rect 1818 6039 1824 6091
rect 1760 5842 1824 6039
rect 1760 5790 1766 5842
rect 1818 5790 1824 5842
rect 1760 5593 1824 5790
rect 1760 5541 1766 5593
rect 1818 5541 1824 5593
rect 1760 5344 1824 5541
rect 1760 5292 1766 5344
rect 1818 5292 1824 5344
rect 1760 5100 1824 5292
rect 1760 5048 1766 5100
rect 1818 5048 1824 5100
rect 1760 4937 1824 5048
rect 3418 7336 3482 7342
rect 3418 7284 3424 7336
rect 3476 7284 3482 7336
rect 3418 7087 3482 7284
rect 3418 7035 3424 7087
rect 3476 7035 3482 7087
rect 3418 6838 3482 7035
rect 3418 6786 3424 6838
rect 3476 6786 3482 6838
rect 3418 6589 3482 6786
rect 3418 6537 3424 6589
rect 3476 6537 3482 6589
rect 3418 6340 3482 6537
rect 3418 6288 3424 6340
rect 3476 6288 3482 6340
rect 3418 6091 3482 6288
rect 5076 7336 5140 7458
rect 8392 7510 8456 7516
rect 8392 7458 8398 7510
rect 8450 7458 8456 7510
rect 5076 7284 5082 7336
rect 5134 7284 5140 7336
rect 5076 7087 5140 7284
rect 5076 7035 5082 7087
rect 5134 7035 5140 7087
rect 5076 6838 5140 7035
rect 5076 6786 5082 6838
rect 5134 6786 5140 6838
rect 5076 6589 5140 6786
rect 5076 6537 5082 6589
rect 5134 6537 5140 6589
rect 5076 6340 5140 6537
rect 5076 6288 5082 6340
rect 5134 6288 5140 6340
rect 3418 6039 3424 6091
rect 3476 6039 3482 6091
rect 3418 5842 3482 6039
rect 3418 5790 3424 5842
rect 3476 5790 3482 5842
rect 3418 5593 3482 5790
rect 3418 5541 3424 5593
rect 3476 5541 3482 5593
rect 3418 5344 3482 5541
rect 3418 5292 3424 5344
rect 3476 5292 3482 5344
rect 3418 5075 3482 5292
rect 4300 6234 4364 6240
rect 4300 6182 4306 6234
rect 4358 6182 4364 6234
rect 4300 5985 4364 6182
rect 4300 5933 4306 5985
rect 4358 5933 4364 5985
rect 4300 5736 4364 5933
rect 4300 5684 4306 5736
rect 4358 5684 4364 5736
rect 4300 5487 4364 5684
rect 4300 5435 4306 5487
rect 4358 5435 4364 5487
rect 4300 5238 4364 5435
rect 4300 5186 4306 5238
rect 4358 5186 4364 5238
rect 3418 5011 3678 5075
rect 1760 4885 1766 4937
rect 1818 4885 1824 4937
rect 1760 4879 1824 4885
rect 3418 4807 3482 4813
rect 3418 4755 3424 4807
rect 3476 4755 3482 4807
rect 3418 4749 3482 4755
rect -1831 4689 -1767 4695
rect -1831 4637 -1825 4689
rect -1773 4637 -1767 4689
rect -1831 4458 -1767 4637
rect -1831 4406 -1825 4458
rect -1773 4406 -1767 4458
rect -1831 4102 -1767 4406
rect 97 4338 171 4347
rect 97 4282 106 4338
rect 162 4282 171 4338
rect 97 4273 171 4282
rect -1831 4050 -1825 4102
rect -1773 4050 -1767 4102
rect -1831 3809 -1767 4050
rect -1831 3757 -1825 3809
rect -1773 3757 -1767 3809
rect -1831 3751 -1767 3757
rect 102 4177 166 4273
rect 102 4125 108 4177
rect 160 4125 166 4177
rect 102 3946 166 4125
rect 102 3894 108 3946
rect 160 3894 166 3946
rect 102 3590 166 3894
rect 102 3538 108 3590
rect 160 3538 166 3590
rect 102 3297 166 3538
rect 102 3245 108 3297
rect 160 3245 166 3297
rect 102 1879 166 3245
rect 1760 4177 1824 4183
rect 1760 4125 1766 4177
rect 1818 4125 1824 4177
rect 1760 3946 1824 4125
rect 3424 3952 3476 4749
rect 1760 3894 1766 3946
rect 1818 3894 1824 3946
rect 1760 3590 1824 3894
rect 3418 3946 3482 3952
rect 3418 3894 3424 3946
rect 3476 3894 3482 3946
rect 3418 3888 3482 3894
rect 1760 3538 1766 3590
rect 1818 3538 1824 3590
rect 1760 3297 1824 3538
rect 3418 3590 3482 3596
rect 3418 3538 3424 3590
rect 3476 3538 3482 3590
rect 3418 3532 3482 3538
rect 1760 3245 1766 3297
rect 1818 3245 1824 3297
rect 1760 3239 1824 3245
rect 3133 2915 3207 2924
rect 3133 2859 3142 2915
rect 3198 2859 3207 2915
rect 3133 2850 3207 2859
rect 1755 2315 1829 2324
rect 1755 2259 1764 2315
rect 1820 2259 1829 2315
rect 1755 2250 1829 2259
rect 102 1827 108 1879
rect 160 1827 166 1879
rect 102 1639 166 1827
rect 1766 1879 1818 2250
rect 3144 1982 3196 2850
rect 3614 2724 3678 5011
rect 4300 4705 4364 5186
rect 5076 6091 5140 6288
rect 6734 7336 6798 7342
rect 6734 7284 6740 7336
rect 6792 7284 6798 7336
rect 6734 7087 6798 7284
rect 6734 7035 6740 7087
rect 6792 7035 6798 7087
rect 6734 6838 6798 7035
rect 6734 6786 6740 6838
rect 6792 6786 6798 6838
rect 6734 6589 6798 6786
rect 6734 6537 6740 6589
rect 6792 6537 6798 6589
rect 6734 6340 6798 6537
rect 6734 6288 6740 6340
rect 6792 6288 6798 6340
rect 5076 6039 5082 6091
rect 5134 6039 5140 6091
rect 5076 5842 5140 6039
rect 5076 5790 5082 5842
rect 5134 5790 5140 5842
rect 5076 5593 5140 5790
rect 5076 5541 5082 5593
rect 5134 5541 5140 5593
rect 5076 5344 5140 5541
rect 5076 5292 5082 5344
rect 5134 5292 5140 5344
rect 5076 5100 5140 5292
rect 5076 5048 5082 5100
rect 5134 5048 5140 5100
rect 5076 4937 5140 5048
rect 5076 4885 5082 4937
rect 5134 4885 5140 4937
rect 5076 4879 5140 4885
rect 5956 6234 6020 6240
rect 5956 6182 5962 6234
rect 6014 6182 6020 6234
rect 5956 5985 6020 6182
rect 5956 5933 5962 5985
rect 6014 5933 6020 5985
rect 5956 5736 6020 5933
rect 5956 5684 5962 5736
rect 6014 5684 6020 5736
rect 5956 5487 6020 5684
rect 5956 5435 5962 5487
rect 6014 5435 6020 5487
rect 5956 5238 6020 5435
rect 5956 5186 5962 5238
rect 6014 5186 6020 5238
rect 4300 4653 4306 4705
rect 4358 4653 4364 4705
rect 3609 2715 3683 2724
rect 3609 2659 3618 2715
rect 3674 2659 3683 2715
rect 3609 2650 3683 2659
rect 3413 2515 3487 2524
rect 3413 2459 3422 2515
rect 3478 2459 3487 2515
rect 3413 2450 3487 2459
rect 3424 2120 3476 2450
rect 4300 2324 4364 4653
rect 5956 4705 6020 5186
rect 6734 6091 6798 6288
rect 6734 6039 6740 6091
rect 6792 6039 6798 6091
rect 6734 5842 6798 6039
rect 6734 5790 6740 5842
rect 6792 5790 6798 5842
rect 6734 5593 6798 5790
rect 6734 5541 6740 5593
rect 6792 5541 6798 5593
rect 6734 5344 6798 5541
rect 6734 5292 6740 5344
rect 6792 5292 6798 5344
rect 6734 5075 6798 5292
rect 5956 4653 5962 4705
rect 6014 4653 6020 4705
rect 5071 4338 5145 4347
rect 5071 4282 5080 4338
rect 5136 4282 5145 4338
rect 5071 4273 5145 4282
rect 5076 4177 5140 4273
rect 5076 4125 5082 4177
rect 5134 4125 5140 4177
rect 5076 3946 5140 4125
rect 5076 3894 5082 3946
rect 5134 3894 5140 3946
rect 5076 3590 5140 3894
rect 5076 3538 5082 3590
rect 5134 3538 5140 3590
rect 5076 3297 5140 3538
rect 5076 3245 5082 3297
rect 5134 3245 5140 3297
rect 5076 3239 5140 3245
rect 4720 3115 4794 3124
rect 4720 3059 4729 3115
rect 4785 3059 4794 3115
rect 4720 3050 4794 3059
rect 4295 2315 4369 2324
rect 4295 2259 4304 2315
rect 4360 2259 4369 2315
rect 4295 2250 4369 2259
rect 3418 2114 3482 2120
rect 3418 2062 3424 2114
rect 3476 2062 3482 2114
rect 3418 2056 3482 2062
rect 3138 1976 3202 1982
rect 3138 1924 3144 1976
rect 3196 1924 3202 1976
rect 3138 1918 3202 1924
rect 1766 1821 1818 1827
rect 3144 1742 3196 1918
rect 3424 1879 3476 2056
rect 4731 1982 4783 3050
rect 5071 2715 5145 2724
rect 5956 2721 6020 4653
rect 6538 5011 6798 5075
rect 8392 7336 8456 7458
rect 8392 7284 8398 7336
rect 8450 7284 8456 7336
rect 8392 7087 8456 7284
rect 8392 7035 8398 7087
rect 8450 7035 8456 7087
rect 8392 6838 8456 7035
rect 8392 6786 8398 6838
rect 8450 6786 8456 6838
rect 8392 6589 8456 6786
rect 8392 6537 8398 6589
rect 8450 6537 8456 6589
rect 8392 6340 8456 6537
rect 8392 6288 8398 6340
rect 8450 6288 8456 6340
rect 8392 6091 8456 6288
rect 8392 6039 8398 6091
rect 8450 6039 8456 6091
rect 8392 5842 8456 6039
rect 8392 5790 8398 5842
rect 8450 5790 8456 5842
rect 8392 5593 8456 5790
rect 8392 5541 8398 5593
rect 8450 5541 8456 5593
rect 8392 5344 8456 5541
rect 8392 5292 8398 5344
rect 8450 5292 8456 5344
rect 8392 5100 8456 5292
rect 8392 5048 8398 5100
rect 8450 5048 8456 5100
rect 5071 2659 5080 2715
rect 5136 2659 5145 2715
rect 5071 2650 5145 2659
rect 5950 2712 6024 2721
rect 5950 2656 5959 2712
rect 6015 2656 6024 2712
rect 4725 1976 4789 1982
rect 4725 1924 4731 1976
rect 4783 1924 4789 1976
rect 4725 1918 4789 1924
rect 3424 1821 3476 1827
rect 4731 1742 4783 1918
rect 5082 1879 5134 2650
rect 5950 2647 6024 2656
rect 6538 2324 6602 5011
rect 8392 4937 8456 5048
rect 8392 4885 8398 4937
rect 8450 4885 8456 4937
rect 8392 4879 8456 4885
rect 10050 7510 10114 7516
rect 10050 7458 10056 7510
rect 10108 7458 10114 7510
rect 10050 7336 10114 7458
rect 10050 7284 10056 7336
rect 10108 7284 10114 7336
rect 10050 7087 10114 7284
rect 10050 7035 10056 7087
rect 10108 7035 10114 7087
rect 10050 6838 10114 7035
rect 10050 6786 10056 6838
rect 10108 6786 10114 6838
rect 10050 6589 10114 6786
rect 10050 6537 10056 6589
rect 10108 6537 10114 6589
rect 10050 6340 10114 6537
rect 10050 6288 10056 6340
rect 10108 6288 10114 6340
rect 10050 6091 10114 6288
rect 10050 6039 10056 6091
rect 10108 6039 10114 6091
rect 10050 5842 10114 6039
rect 10050 5790 10056 5842
rect 10108 5790 10114 5842
rect 10050 5593 10114 5790
rect 10050 5541 10056 5593
rect 10108 5541 10114 5593
rect 10050 5344 10114 5541
rect 10050 5292 10056 5344
rect 10108 5292 10114 5344
rect 10050 5100 10114 5292
rect 10050 5048 10056 5100
rect 10108 5048 10114 5100
rect 10050 4937 10114 5048
rect 10050 4885 10056 4937
rect 10108 4885 10114 4937
rect 10050 4879 10114 4885
rect 6734 4807 6798 4813
rect 6734 4755 6740 4807
rect 6792 4755 6798 4807
rect 6734 4749 6798 4755
rect 6740 3952 6792 4749
rect 10045 4338 10119 4347
rect 10045 4282 10054 4338
rect 10110 4282 10119 4338
rect 10045 4273 10119 4282
rect 8392 4177 8456 4183
rect 8392 4125 8398 4177
rect 8450 4125 8456 4177
rect 6734 3946 6798 3952
rect 6734 3894 6740 3946
rect 6792 3894 6798 3946
rect 6734 3888 6798 3894
rect 8392 3946 8456 4125
rect 8392 3894 8398 3946
rect 8450 3894 8456 3946
rect 8392 3590 8456 3894
rect 8392 3538 8398 3590
rect 8450 3538 8456 3590
rect 6734 3466 6798 3472
rect 6734 3414 6740 3466
rect 6792 3414 6798 3466
rect 6734 3408 6798 3414
rect 6740 2524 6792 3408
rect 8392 3297 8456 3538
rect 8392 3245 8398 3297
rect 8450 3245 8456 3297
rect 8392 3239 8456 3245
rect 10050 4177 10114 4273
rect 10050 4125 10056 4177
rect 10108 4125 10114 4177
rect 10050 3946 10114 4125
rect 10050 3894 10056 3946
rect 10108 3894 10114 3946
rect 10050 3590 10114 3894
rect 10050 3538 10056 3590
rect 10108 3538 10114 3590
rect 10050 3297 10114 3538
rect 10050 3245 10056 3297
rect 10108 3245 10114 3297
rect 6952 2915 7026 2924
rect 6952 2859 6961 2915
rect 7017 2859 7026 2915
rect 6952 2850 7026 2859
rect 6729 2515 6803 2524
rect 6729 2459 6738 2515
rect 6794 2459 6803 2515
rect 6729 2450 6803 2459
rect 6533 2315 6607 2324
rect 6533 2259 6542 2315
rect 6598 2259 6607 2315
rect 6533 2250 6607 2259
rect 6740 2120 6792 2450
rect 6734 2114 6798 2120
rect 6734 2062 6740 2114
rect 6792 2062 6798 2114
rect 6734 2056 6798 2062
rect 5082 1821 5134 1827
rect 6740 1879 6792 2056
rect 6963 1982 7015 2850
rect 8387 2315 8461 2324
rect 8387 2259 8396 2315
rect 8452 2259 8461 2315
rect 8387 2250 8461 2259
rect 6957 1976 7021 1982
rect 6957 1924 6963 1976
rect 7015 1924 7021 1976
rect 6957 1918 7021 1924
rect 6740 1821 6792 1827
rect 6963 1742 7015 1918
rect 8398 1879 8450 2250
rect 8398 1821 8450 1827
rect 10050 1879 10114 3245
rect 10050 1827 10056 1879
rect 10108 1827 10114 1879
rect 3138 1736 3202 1742
rect 3138 1684 3144 1736
rect 3196 1684 3202 1736
rect 3138 1678 3202 1684
rect 4725 1736 4789 1742
rect 4725 1684 4731 1736
rect 4783 1684 4789 1736
rect 4725 1678 4789 1684
rect 6957 1736 7021 1742
rect 6957 1684 6963 1736
rect 7015 1684 7021 1736
rect 6957 1678 7021 1684
rect 102 1587 108 1639
rect 160 1587 166 1639
rect 102 1399 166 1587
rect 1766 1639 1818 1645
rect 1766 1581 1818 1587
rect 3144 1502 3196 1678
rect 3424 1639 3476 1645
rect 3424 1581 3476 1587
rect 4731 1502 4783 1678
rect 5082 1639 5134 1645
rect 5082 1581 5134 1587
rect 6740 1639 6792 1645
rect 6740 1581 6792 1587
rect 6963 1502 7015 1678
rect 8398 1639 8450 1645
rect 8398 1581 8450 1587
rect 10050 1639 10114 1827
rect 10050 1587 10056 1639
rect 10108 1587 10114 1639
rect 3138 1496 3202 1502
rect 3138 1444 3144 1496
rect 3196 1444 3202 1496
rect 3138 1438 3202 1444
rect 4725 1496 4789 1502
rect 4725 1444 4731 1496
rect 4783 1444 4789 1496
rect 4725 1438 4789 1444
rect 6957 1496 7021 1502
rect 6957 1444 6963 1496
rect 7015 1444 7021 1496
rect 6957 1438 7021 1444
rect 102 1347 108 1399
rect 160 1347 166 1399
rect 102 1159 166 1347
rect 1766 1399 1818 1405
rect 1766 1341 1818 1347
rect 3144 1262 3196 1438
rect 3424 1399 3476 1405
rect 3424 1341 3476 1347
rect 4731 1262 4783 1438
rect 5082 1399 5134 1405
rect 5082 1341 5134 1347
rect 6740 1399 6792 1405
rect 6740 1341 6792 1347
rect 6963 1262 7015 1438
rect 8398 1399 8450 1405
rect 8398 1341 8450 1347
rect 10050 1399 10114 1587
rect 10050 1347 10056 1399
rect 10108 1347 10114 1399
rect 3138 1256 3202 1262
rect 3138 1204 3144 1256
rect 3196 1204 3202 1256
rect 3138 1198 3202 1204
rect 4725 1256 4789 1262
rect 4725 1204 4731 1256
rect 4783 1204 4789 1256
rect 4725 1198 4789 1204
rect 6957 1256 7021 1262
rect 6957 1204 6963 1256
rect 7015 1204 7021 1256
rect 6957 1198 7021 1204
rect 102 1107 108 1159
rect 160 1107 166 1159
rect 102 919 166 1107
rect 1766 1159 1818 1165
rect 1766 1101 1818 1107
rect 3144 1022 3196 1198
rect 3424 1159 3476 1165
rect 3424 1101 3476 1107
rect 4731 1022 4783 1198
rect 5082 1159 5134 1165
rect 5082 1101 5134 1107
rect 6740 1159 6792 1165
rect 6740 1101 6792 1107
rect 6963 1022 7015 1198
rect 8398 1159 8450 1165
rect 8398 1101 8450 1107
rect 10050 1159 10114 1347
rect 10050 1107 10056 1159
rect 10108 1107 10114 1159
rect 3138 1016 3202 1022
rect 3138 964 3144 1016
rect 3196 964 3202 1016
rect 3138 958 3202 964
rect 4725 1016 4789 1022
rect 4725 964 4731 1016
rect 4783 964 4789 1016
rect 4725 958 4789 964
rect 6957 1016 7021 1022
rect 6957 964 6963 1016
rect 7015 964 7021 1016
rect 6957 958 7021 964
rect 102 867 108 919
rect 160 867 166 919
rect 102 679 166 867
rect 1766 919 1818 925
rect 1766 861 1818 867
rect 3144 782 3196 958
rect 3424 919 3476 925
rect 3424 861 3476 867
rect 4731 782 4783 958
rect 5082 919 5134 925
rect 5082 861 5134 867
rect 6740 919 6792 925
rect 6740 861 6792 867
rect 6963 782 7015 958
rect 8398 919 8450 925
rect 8398 861 8450 867
rect 10050 919 10114 1107
rect 10050 867 10056 919
rect 10108 867 10114 919
rect 3138 776 3202 782
rect 3138 724 3144 776
rect 3196 724 3202 776
rect 3138 718 3202 724
rect 4725 776 4789 782
rect 4725 724 4731 776
rect 4783 724 4789 776
rect 4725 718 4789 724
rect 6957 776 7021 782
rect 6957 724 6963 776
rect 7015 724 7021 776
rect 6957 718 7021 724
rect 102 627 108 679
rect 160 627 166 679
rect 102 439 166 627
rect 1766 679 1818 685
rect 1766 621 1818 627
rect 3144 542 3196 718
rect 3424 679 3476 685
rect 3424 621 3476 627
rect 4731 542 4783 718
rect 5082 679 5134 685
rect 5082 621 5134 627
rect 6740 679 6792 685
rect 6740 621 6792 627
rect 6963 542 7015 718
rect 8398 679 8450 685
rect 8398 621 8450 627
rect 10050 679 10114 867
rect 10050 627 10056 679
rect 10108 627 10114 679
rect 3138 536 3202 542
rect 3138 484 3144 536
rect 3196 484 3202 536
rect 3138 478 3202 484
rect 4725 536 4789 542
rect 4725 484 4731 536
rect 4783 484 4789 536
rect 4725 478 4789 484
rect 6957 536 7021 542
rect 6957 484 6963 536
rect 7015 484 7021 536
rect 6957 478 7021 484
rect 102 387 108 439
rect 160 387 166 439
rect 102 199 166 387
rect 1766 439 1818 445
rect 1766 381 1818 387
rect 3144 302 3196 478
rect 3424 439 3476 445
rect 3424 381 3476 387
rect 4731 302 4783 478
rect 5082 439 5134 445
rect 5082 381 5134 387
rect 6740 439 6792 445
rect 6740 381 6792 387
rect 6963 302 7015 478
rect 8398 439 8450 445
rect 8398 381 8450 387
rect 10050 439 10114 627
rect 10050 387 10056 439
rect 10108 387 10114 439
rect 3138 296 3202 302
rect 3138 244 3144 296
rect 3196 244 3202 296
rect 3138 238 3202 244
rect 4725 296 4789 302
rect 4725 244 4731 296
rect 4783 244 4789 296
rect 4725 238 4789 244
rect 6957 296 7021 302
rect 6957 244 6963 296
rect 7015 244 7021 296
rect 6957 238 7021 244
rect 102 147 108 199
rect 160 147 166 199
rect 102 -77 166 147
rect 1766 199 1818 205
rect 1766 141 1818 147
rect 3424 199 3476 205
rect 3424 32 3476 147
rect 5082 199 5134 205
rect 5082 141 5134 147
rect 6740 199 6792 205
rect 3418 26 3482 32
rect 6740 31 6792 147
rect 8398 199 8450 205
rect 8398 141 8450 147
rect 10050 199 10114 387
rect 10050 147 10056 199
rect 10108 147 10114 199
rect 3418 -26 3424 26
rect 3476 -26 3482 26
rect 3418 -32 3482 -26
rect 6734 25 6798 31
rect 6734 -27 6740 25
rect 6792 -27 6798 25
rect 6734 -33 6798 -27
rect 10050 -77 10114 147
rect 97 -86 171 -77
rect 97 -142 106 -86
rect 162 -142 171 -86
rect 97 -151 171 -142
rect 10045 -86 10119 -77
rect 10045 -142 10054 -86
rect 10110 -142 10119 -86
rect 10045 -151 10119 -142
<< via2 >>
rect -1030 6196 -974 6252
rect 106 4282 162 4338
rect 3142 2859 3198 2915
rect 1764 2259 1820 2315
rect 3618 2659 3674 2715
rect 3422 2459 3478 2515
rect 5080 4282 5136 4338
rect 4729 3059 4785 3115
rect 4304 2259 4360 2315
rect 5080 2659 5136 2715
rect 5959 2656 6015 2712
rect 10054 4282 10110 4338
rect 6961 2859 7017 2915
rect 6738 2459 6794 2515
rect 6542 2259 6598 2315
rect 8396 2259 8452 2315
rect 106 -142 162 -86
rect 10054 -142 10110 -86
<< metal3 >>
rect -1039 6252 -965 6261
rect -1039 6196 -1030 6252
rect -974 6196 -965 6252
rect -1039 6187 -965 6196
rect 97 4340 171 4347
rect 5071 4340 5145 4347
rect 10045 4340 10119 4347
rect 97 4338 10119 4340
rect 97 4282 106 4338
rect 162 4282 5080 4338
rect 5136 4282 10054 4338
rect 10110 4282 10119 4338
rect 97 4280 10119 4282
rect 97 4273 171 4280
rect 5071 4273 5145 4280
rect 10045 4273 10119 4280
rect 4720 3117 4794 3124
rect 1766 3115 8450 3117
rect 1766 3059 4729 3115
rect 4785 3059 8450 3115
rect 1766 3057 8450 3059
rect 4720 3050 4794 3057
rect 3133 2917 3207 2924
rect 6952 2917 7026 2924
rect 1766 2915 8450 2917
rect 1766 2859 3142 2915
rect 3198 2859 6961 2915
rect 7017 2859 8450 2915
rect 1766 2857 8450 2859
rect 3133 2850 3207 2857
rect 6952 2850 7026 2857
rect 3609 2717 3683 2724
rect 5071 2717 5145 2724
rect 5950 2717 6024 2721
rect 1766 2715 8450 2717
rect 1766 2659 3618 2715
rect 3674 2659 5080 2715
rect 5136 2712 8450 2715
rect 5136 2659 5959 2712
rect 1766 2657 5959 2659
rect 3609 2650 3683 2657
rect 5071 2650 5145 2657
rect 5950 2656 5959 2657
rect 6015 2657 8450 2712
rect 6015 2656 6024 2657
rect 5950 2647 6024 2656
rect 3413 2517 3487 2524
rect 6729 2517 6803 2524
rect 1766 2515 8450 2517
rect 1766 2459 3422 2515
rect 3478 2459 6738 2515
rect 6794 2459 8450 2515
rect 1766 2457 8450 2459
rect 3413 2450 3487 2457
rect 6729 2450 6803 2457
rect 1755 2317 1829 2324
rect 4295 2317 4369 2324
rect 6533 2317 6607 2324
rect 8387 2317 8461 2324
rect 1755 2315 8461 2317
rect 1755 2259 1764 2315
rect 1820 2259 4304 2315
rect 4360 2259 6542 2315
rect 6598 2259 8396 2315
rect 8452 2259 8461 2315
rect 1755 2257 8461 2259
rect 1755 2250 1829 2257
rect 4295 2250 4369 2257
rect 6533 2250 6607 2257
rect 8387 2250 8461 2257
rect 97 -84 171 -77
rect 10045 -84 10119 -77
rect 97 -86 10119 -84
rect 97 -142 106 -86
rect 162 -142 10054 -86
rect 10110 -142 10119 -86
rect 97 -144 10119 -142
rect 97 -151 171 -144
rect 10045 -151 10119 -144
use sky130_fd_pr__nfet_g5v0d10v5_GLAJGT  sky130_fd_pr__nfet_g5v0d10v5_GLAJGT_1
timestamp 1711730665
transform 1 0 5108 0 1 1044
box -5173 -1109 5173 1109
use sky130_fd_pr__nfet_g5v0d10v5_T82T27  sky130_fd_pr__nfet_g5v0d10v5_T82T27_1
timestamp 1711813642
transform 1 0 5108 0 1 3711
box -5173 -505 5173 505
use sky130_fd_pr__pfet_g5v0d10v5_3HV7M9  sky130_fd_pr__pfet_g5v0d10v5_3HV7M9_0
timestamp 1711774300
transform 1 0 5108 0 1 4807
box -5203 -362 5203 362
use sky130_fd_pr__pfet_g5v0d10v5_8FRRWQ  sky130_fd_pr__pfet_g5v0d10v5_8FRRWQ_0
timestamp 1711767182
transform 1 0 5108 0 1 6279
box -5203 -1300 5203 1300
<< labels >>
rlabel metal3 1755 2317 1755 2317 7 vnn
rlabel metal3 1766 2717 1766 2717 7 vpp
rlabel metal3 1766 2917 1766 2917 7 vinn
port 1 w
rlabel metal3 1766 3117 1766 3117 7 vinp
port 2 w
rlabel metal3 97 -84 97 -84 7 avss
port 3 w
rlabel metal3 1766 2517 1766 2517 7 vt
rlabel metal2 102 7516 102 7516 7 avdd
port 4 w
rlabel metal2 3424 4230 3424 4230 7 vm
rlabel metal2 6740 4230 6740 4230 7 n0
rlabel metal2 3418 3596 3418 3596 7 vn
<< end >>
