magic
tech sky130A
magscale 1 2
timestamp 1711636687
<< mvnmos >>
rect -60 -73 60 11
<< mvndiff >>
rect -118 -1 -60 11
rect -118 -61 -106 -1
rect -72 -61 -60 -1
rect -118 -73 -60 -61
rect 60 -1 118 11
rect 60 -61 72 -1
rect 106 -61 118 -1
rect 60 -73 118 -61
<< mvndiffc >>
rect -106 -61 -72 -1
rect 72 -61 106 -1
<< poly >>
rect -60 83 60 99
rect -60 49 -44 83
rect 44 49 60 83
rect -60 11 60 49
rect -60 -99 60 -73
<< polycont >>
rect -44 49 44 83
<< locali >>
rect -60 49 -44 83
rect 44 49 60 83
rect -106 -1 -72 15
rect -106 -77 -72 -61
rect 72 -1 106 15
rect 72 -77 106 -61
<< viali >>
rect -44 49 44 83
rect -106 -61 -72 -1
rect 72 -61 106 -1
<< metal1 >>
rect -56 83 56 89
rect -56 49 -44 83
rect 44 49 56 83
rect -56 43 56 49
rect -112 -1 -66 11
rect -112 -61 -106 -1
rect -72 -61 -66 -1
rect -112 -73 -66 -61
rect 66 -1 112 11
rect 66 -61 72 -1
rect 106 -61 112 -1
rect 66 -73 112 -61
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.60 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
