magic
tech sky130A
magscale 1 2
timestamp 1712531369
<< viali >>
rect 1685 7361 1719 7395
rect 10241 7361 10275 7395
rect 1501 7157 1535 7191
rect 10425 7157 10459 7191
rect 2145 6409 2179 6443
rect 2881 6341 2915 6375
rect 1685 6273 1719 6307
rect 10241 6273 10275 6307
rect 2329 6205 2363 6239
rect 2421 6205 2455 6239
rect 9689 6205 9723 6239
rect 9781 6205 9815 6239
rect 9873 6205 9907 6239
rect 9965 6205 9999 6239
rect 1501 6137 1535 6171
rect 2881 6137 2915 6171
rect 10425 6137 10459 6171
rect 9505 6069 9539 6103
rect 1685 5865 1719 5899
rect 10241 5865 10275 5899
rect 2421 5797 2455 5831
rect 3341 5797 3375 5831
rect 1869 5729 1903 5763
rect 9873 5729 9907 5763
rect 10082 5729 10116 5763
rect 2605 5661 2639 5695
rect 9505 5661 9539 5695
rect 9597 5661 9631 5695
rect 9965 5661 9999 5695
rect 2421 5593 2455 5627
rect 2789 5593 2823 5627
rect 3341 5593 3375 5627
rect 1961 5525 1995 5559
rect 2881 5525 2915 5559
rect 9321 5525 9355 5559
rect 1501 5321 1535 5355
rect 9965 5321 9999 5355
rect 10241 5321 10275 5355
rect 1685 5185 1719 5219
rect 2053 5185 2087 5219
rect 9505 5185 9539 5219
rect 10082 5185 10116 5219
rect 9597 5117 9631 5151
rect 9873 5117 9907 5151
rect 1869 4981 1903 5015
rect 9321 4981 9355 5015
rect 2053 4777 2087 4811
rect 9597 4777 9631 4811
rect 2789 4709 2823 4743
rect 10241 4641 10275 4675
rect 1685 4573 1719 4607
rect 9505 4573 9539 4607
rect 9965 4573 9999 4607
rect 2789 4505 2823 4539
rect 9756 4505 9790 4539
rect 1501 4437 1535 4471
rect 2237 4437 2271 4471
rect 2329 4437 2363 4471
rect 9321 4437 9355 4471
rect 9873 4437 9907 4471
rect 2421 4233 2455 4267
rect 2605 4233 2639 4267
rect 9689 4233 9723 4267
rect 9965 4233 9999 4267
rect 10333 4233 10367 4267
rect 3157 4165 3191 4199
rect 2697 4097 2731 4131
rect 9873 4097 9907 4131
rect 10057 4097 10091 4131
rect 10517 4097 10551 4131
rect 3157 3961 3191 3995
rect 10241 3961 10275 3995
rect 9321 3689 9355 3723
rect 10333 3689 10367 3723
rect 9597 3621 9631 3655
rect 9965 3553 9999 3587
rect 10241 3553 10275 3587
rect 6285 3485 6319 3519
rect 9505 3485 9539 3519
rect 9756 3485 9790 3519
rect 10517 3485 10551 3519
rect 6469 3349 6503 3383
rect 9873 3349 9907 3383
rect 5457 3145 5491 3179
rect 5549 3077 5583 3111
rect 6561 3077 6595 3111
rect 6653 3077 6687 3111
rect 7113 3077 7147 3111
rect 9597 3077 9631 3111
rect 10057 3077 10091 3111
rect 3617 3009 3651 3043
rect 3709 3009 3743 3043
rect 4169 3009 4203 3043
rect 4461 3009 4495 3043
rect 4813 3009 4847 3043
rect 5917 3009 5951 3043
rect 9505 3009 9539 3043
rect 10241 3009 10275 3043
rect 3525 2941 3559 2975
rect 3801 2941 3835 2975
rect 4261 2941 4295 2975
rect 4353 2941 4387 2975
rect 4629 2941 4663 2975
rect 4905 2941 4939 2975
rect 4997 2941 5031 2975
rect 5089 2941 5123 2975
rect 9965 2941 9999 2975
rect 5733 2873 5767 2907
rect 7113 2873 7147 2907
rect 9597 2873 9631 2907
rect 9873 2873 9907 2907
rect 3985 2805 4019 2839
rect 5273 2805 5307 2839
rect 6377 2805 6411 2839
rect 9321 2805 9355 2839
rect 9781 2805 9815 2839
rect 6561 2601 6595 2635
rect 7389 2601 7423 2635
rect 8033 2601 8067 2635
rect 8677 2533 8711 2567
rect 9965 2533 9999 2567
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 6193 2397 6227 2431
rect 6377 2397 6411 2431
rect 6837 2397 6871 2431
rect 7205 2397 7239 2431
rect 7849 2397 7883 2431
rect 8493 2397 8527 2431
rect 10149 2397 10183 2431
rect 4169 2261 4203 2295
rect 4813 2261 4847 2295
rect 5457 2261 5491 2295
rect 6009 2261 6043 2295
rect 6653 2261 6687 2295
<< metal1 >>
rect 1104 9818 10856 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 10856 9818
rect 1104 9744 10856 9766
rect 1104 9274 10856 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 10856 9274
rect 1104 9200 10856 9222
rect 1104 8730 10856 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 10856 8730
rect 1104 8656 10856 8678
rect 1104 8186 10856 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 10856 8186
rect 1104 8112 10856 8134
rect 1104 7642 10856 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 10856 7642
rect 1104 7568 10856 7590
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 10226 7352 10232 7404
rect 10284 7352 10290 7404
rect 1486 7148 1492 7200
rect 1544 7148 1550 7200
rect 10410 7148 10416 7200
rect 10468 7148 10474 7200
rect 1104 7098 10856 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 10856 7098
rect 1104 7024 10856 7046
rect 1104 6554 10856 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 10856 6554
rect 1104 6480 10856 6502
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 1728 6412 2145 6440
rect 1728 6400 1734 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 2869 6375 2927 6381
rect 2869 6341 2881 6375
rect 2915 6341 2927 6375
rect 2869 6335 2927 6341
rect 1670 6264 1676 6316
rect 1728 6264 1734 6316
rect 2884 6304 2912 6335
rect 3050 6304 3056 6316
rect 2884 6276 3056 6304
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 10192 6276 10241 6304
rect 10192 6264 10198 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 2314 6196 2320 6248
rect 2372 6196 2378 6248
rect 2406 6196 2412 6248
rect 2464 6196 2470 6248
rect 9674 6196 9680 6248
rect 9732 6196 9738 6248
rect 9766 6196 9772 6248
rect 9824 6196 9830 6248
rect 9861 6239 9919 6245
rect 9861 6205 9873 6239
rect 9907 6205 9919 6239
rect 9861 6199 9919 6205
rect 934 6128 940 6180
rect 992 6168 998 6180
rect 1489 6171 1547 6177
rect 1489 6168 1501 6171
rect 992 6140 1501 6168
rect 992 6128 998 6140
rect 1489 6137 1501 6140
rect 1535 6137 1547 6171
rect 1489 6131 1547 6137
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 2958 6168 2964 6180
rect 2915 6140 2964 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 9876 6168 9904 6199
rect 9950 6196 9956 6248
rect 10008 6196 10014 6248
rect 10042 6196 10048 6248
rect 10100 6196 10106 6248
rect 10060 6168 10088 6196
rect 9876 6140 10088 6168
rect 10410 6128 10416 6180
rect 10468 6128 10474 6180
rect 9490 6060 9496 6112
rect 9548 6060 9554 6112
rect 1104 6010 10856 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 10856 6010
rect 1104 5936 10856 5958
rect 1670 5856 1676 5908
rect 1728 5856 1734 5908
rect 9490 5856 9496 5908
rect 9548 5856 9554 5908
rect 9858 5856 9864 5908
rect 9916 5856 9922 5908
rect 10226 5856 10232 5908
rect 10284 5856 10290 5908
rect 2314 5788 2320 5840
rect 2372 5828 2378 5840
rect 2409 5831 2467 5837
rect 2409 5828 2421 5831
rect 2372 5800 2421 5828
rect 2372 5788 2378 5800
rect 2409 5797 2421 5800
rect 2455 5828 2467 5831
rect 2774 5828 2780 5840
rect 2455 5800 2780 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 2774 5788 2780 5800
rect 2832 5788 2838 5840
rect 2958 5828 2964 5840
rect 2884 5800 2964 5828
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 2884 5760 2912 5800
rect 2958 5788 2964 5800
rect 3016 5828 3022 5840
rect 3329 5831 3387 5837
rect 3329 5828 3341 5831
rect 3016 5800 3341 5828
rect 3016 5788 3022 5800
rect 3329 5797 3341 5800
rect 3375 5797 3387 5831
rect 3329 5791 3387 5797
rect 1903 5732 2912 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 9508 5701 9536 5856
rect 9876 5828 9904 5856
rect 9876 5800 9996 5828
rect 9674 5720 9680 5772
rect 9732 5720 9738 5772
rect 9766 5720 9772 5772
rect 9824 5760 9830 5772
rect 9861 5763 9919 5769
rect 9861 5760 9873 5763
rect 9824 5732 9873 5760
rect 9824 5720 9830 5732
rect 9861 5729 9873 5732
rect 9907 5729 9919 5763
rect 9968 5760 9996 5800
rect 10070 5763 10128 5769
rect 10070 5760 10082 5763
rect 9968 5732 10082 5760
rect 9861 5723 9919 5729
rect 10070 5729 10082 5732
rect 10116 5729 10128 5763
rect 10070 5723 10128 5729
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 1820 5664 2605 5692
rect 1820 5652 1826 5664
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 9585 5695 9643 5701
rect 9585 5661 9597 5695
rect 9631 5661 9643 5695
rect 9692 5692 9720 5720
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9692 5664 9965 5692
rect 9585 5655 9643 5661
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 2314 5584 2320 5636
rect 2372 5624 2378 5636
rect 2409 5627 2467 5633
rect 2409 5624 2421 5627
rect 2372 5596 2421 5624
rect 2372 5584 2378 5596
rect 2409 5593 2421 5596
rect 2455 5593 2467 5627
rect 2409 5587 2467 5593
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 3329 5627 3387 5633
rect 2832 5596 3188 5624
rect 2832 5584 2838 5596
rect 3160 5568 3188 5596
rect 3329 5593 3341 5627
rect 3375 5624 3387 5627
rect 3510 5624 3516 5636
rect 3375 5596 3516 5624
rect 3375 5593 3387 5596
rect 3329 5587 3387 5593
rect 3510 5584 3516 5596
rect 3568 5584 3574 5636
rect 9600 5624 9628 5655
rect 9600 5596 10088 5624
rect 10060 5568 10088 5596
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 2869 5559 2927 5565
rect 2869 5556 2881 5559
rect 1995 5528 2881 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 2869 5525 2881 5528
rect 2915 5556 2927 5559
rect 3050 5556 3056 5568
rect 2915 5528 3056 5556
rect 2915 5525 2927 5528
rect 2869 5519 2927 5525
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 3142 5516 3148 5568
rect 3200 5516 3206 5568
rect 9306 5516 9312 5568
rect 9364 5516 9370 5568
rect 10042 5516 10048 5568
rect 10100 5516 10106 5568
rect 1104 5466 10856 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 10856 5466
rect 1104 5392 10856 5414
rect 842 5312 848 5364
rect 900 5352 906 5364
rect 1489 5355 1547 5361
rect 1489 5352 1501 5355
rect 900 5324 1501 5352
rect 900 5312 906 5324
rect 1489 5321 1501 5324
rect 1535 5321 1547 5355
rect 1489 5315 1547 5321
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 9824 5324 9965 5352
rect 9824 5312 9830 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 9953 5315 10011 5321
rect 10134 5312 10140 5364
rect 10192 5352 10198 5364
rect 10229 5355 10287 5361
rect 10229 5352 10241 5355
rect 10192 5324 10241 5352
rect 10192 5312 10198 5324
rect 10229 5321 10241 5324
rect 10275 5321 10287 5355
rect 10229 5315 10287 5321
rect 9674 5244 9680 5296
rect 9732 5244 9738 5296
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 1762 5216 1768 5228
rect 1719 5188 1768 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 1854 5176 1860 5228
rect 1912 5216 1918 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 1912 5188 2053 5216
rect 1912 5176 1918 5188
rect 2041 5185 2053 5188
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 9490 5176 9496 5228
rect 9548 5176 9554 5228
rect 9692 5216 9720 5244
rect 9950 5216 9956 5228
rect 9692 5188 9956 5216
rect 9950 5176 9956 5188
rect 10008 5216 10014 5228
rect 10070 5219 10128 5225
rect 10070 5216 10082 5219
rect 10008 5188 10082 5216
rect 10008 5176 10014 5188
rect 10070 5185 10082 5188
rect 10116 5185 10128 5219
rect 10070 5179 10128 5185
rect 9582 5108 9588 5160
rect 9640 5108 9646 5160
rect 9861 5151 9919 5157
rect 9861 5117 9873 5151
rect 9907 5148 9919 5151
rect 10226 5148 10232 5160
rect 9907 5120 10232 5148
rect 9907 5117 9919 5120
rect 9861 5111 9919 5117
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 992 4984 1869 5012
rect 992 4972 998 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 9306 4972 9312 5024
rect 9364 4972 9370 5024
rect 1104 4922 10856 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 10856 4922
rect 1104 4848 10856 4870
rect 1854 4768 1860 4820
rect 1912 4808 1918 4820
rect 2041 4811 2099 4817
rect 2041 4808 2053 4811
rect 1912 4780 2053 4808
rect 1912 4768 1918 4780
rect 2041 4777 2053 4780
rect 2087 4777 2099 4811
rect 2041 4771 2099 4777
rect 9490 4768 9496 4820
rect 9548 4808 9554 4820
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 9548 4780 9597 4808
rect 9548 4768 9554 4780
rect 9585 4777 9597 4780
rect 9631 4777 9643 4811
rect 9585 4771 9643 4777
rect 2777 4743 2835 4749
rect 2777 4709 2789 4743
rect 2823 4740 2835 4743
rect 3142 4740 3148 4752
rect 2823 4712 3148 4740
rect 2823 4709 2835 4712
rect 2777 4703 2835 4709
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 9674 4672 9680 4684
rect 9508 4644 9680 4672
rect 1670 4564 1676 4616
rect 1728 4564 1734 4616
rect 9508 4613 9536 4644
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 10229 4675 10287 4681
rect 10229 4672 10241 4675
rect 9824 4644 10241 4672
rect 9824 4632 9830 4644
rect 10229 4641 10241 4644
rect 10275 4641 10287 4675
rect 10229 4635 10287 4641
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 9950 4564 9956 4616
rect 10008 4564 10014 4616
rect 2777 4539 2835 4545
rect 2777 4505 2789 4539
rect 2823 4536 2835 4539
rect 2958 4536 2964 4548
rect 2823 4508 2964 4536
rect 2823 4505 2835 4508
rect 2777 4499 2835 4505
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 9744 4539 9802 4545
rect 9744 4505 9756 4539
rect 9790 4536 9802 4539
rect 10042 4536 10048 4548
rect 9790 4508 10048 4536
rect 9790 4505 9802 4508
rect 9744 4499 9802 4505
rect 10042 4496 10048 4508
rect 10100 4496 10106 4548
rect 1486 4428 1492 4480
rect 1544 4428 1550 4480
rect 2222 4428 2228 4480
rect 2280 4428 2286 4480
rect 2314 4428 2320 4480
rect 2372 4428 2378 4480
rect 9306 4428 9312 4480
rect 9364 4428 9370 4480
rect 9858 4428 9864 4480
rect 9916 4428 9922 4480
rect 1104 4378 10856 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 10856 4378
rect 1104 4304 10856 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 2409 4267 2467 4273
rect 2409 4264 2421 4267
rect 1728 4236 2421 4264
rect 1728 4224 1734 4236
rect 2409 4233 2421 4236
rect 2455 4233 2467 4267
rect 2409 4227 2467 4233
rect 2593 4267 2651 4273
rect 2593 4233 2605 4267
rect 2639 4264 2651 4267
rect 2958 4264 2964 4276
rect 2639 4236 2964 4264
rect 2639 4233 2651 4236
rect 2593 4227 2651 4233
rect 2958 4224 2964 4236
rect 3016 4264 3022 4276
rect 3694 4264 3700 4276
rect 3016 4236 3700 4264
rect 3016 4224 3022 4236
rect 3694 4224 3700 4236
rect 3752 4224 3758 4276
rect 9674 4224 9680 4276
rect 9732 4224 9738 4276
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 9953 4267 10011 4273
rect 9953 4264 9965 4267
rect 9824 4236 9965 4264
rect 9824 4224 9830 4236
rect 9953 4233 9965 4236
rect 9999 4264 10011 4267
rect 10321 4267 10379 4273
rect 10321 4264 10333 4267
rect 9999 4236 10333 4264
rect 9999 4233 10011 4236
rect 9953 4227 10011 4233
rect 10321 4233 10333 4236
rect 10367 4233 10379 4267
rect 10321 4227 10379 4233
rect 2222 4156 2228 4208
rect 2280 4196 2286 4208
rect 3050 4196 3056 4208
rect 2280 4168 3056 4196
rect 2280 4156 2286 4168
rect 3050 4156 3056 4168
rect 3108 4196 3114 4208
rect 3145 4199 3203 4205
rect 3145 4196 3157 4199
rect 3108 4168 3157 4196
rect 3108 4156 3114 4168
rect 3145 4165 3157 4168
rect 3191 4196 3203 4199
rect 3191 4168 3924 4196
rect 3191 4165 3203 4168
rect 3145 4159 3203 4165
rect 2314 4088 2320 4140
rect 2372 4128 2378 4140
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2372 4100 2697 4128
rect 2372 4088 2378 4100
rect 2685 4097 2697 4100
rect 2731 4128 2743 4131
rect 2731 4100 3556 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 3528 4072 3556 4100
rect 3896 4072 3924 4168
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 9950 4128 9956 4140
rect 9907 4100 9956 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 10042 4088 10048 4140
rect 10100 4088 10106 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 3510 4020 3516 4072
rect 3568 4020 3574 4072
rect 3878 4020 3884 4072
rect 3936 4020 3942 4072
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 10520 4060 10548 4091
rect 7432 4032 10548 4060
rect 7432 4020 7438 4032
rect 3142 3952 3148 4004
rect 3200 3952 3206 4004
rect 6638 3952 6644 4004
rect 6696 3992 6702 4004
rect 9858 3992 9864 4004
rect 6696 3964 9864 3992
rect 6696 3952 6702 3964
rect 9858 3952 9864 3964
rect 9916 3992 9922 4004
rect 10229 3995 10287 4001
rect 10229 3992 10241 3995
rect 9916 3964 10241 3992
rect 9916 3952 9922 3964
rect 10229 3961 10241 3964
rect 10275 3961 10287 3995
rect 10229 3955 10287 3961
rect 3160 3924 3188 3952
rect 3602 3924 3608 3936
rect 3160 3896 3608 3924
rect 3602 3884 3608 3896
rect 3660 3924 3666 3936
rect 4246 3924 4252 3936
rect 3660 3896 4252 3924
rect 3660 3884 3666 3896
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 1104 3834 10856 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 10856 3834
rect 1104 3760 10856 3782
rect 9309 3723 9367 3729
rect 9309 3689 9321 3723
rect 9355 3689 9367 3723
rect 9309 3683 9367 3689
rect 9324 3596 9352 3683
rect 9766 3680 9772 3732
rect 9824 3680 9830 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10321 3723 10379 3729
rect 10321 3720 10333 3723
rect 10008 3692 10333 3720
rect 10008 3680 10014 3692
rect 9585 3655 9643 3661
rect 9585 3621 9597 3655
rect 9631 3621 9643 3655
rect 9585 3615 9643 3621
rect 9306 3544 9312 3596
rect 9364 3544 9370 3596
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3516 6331 3519
rect 9493 3519 9551 3525
rect 6319 3488 6408 3516
rect 6319 3485 6331 3488
rect 6273 3479 6331 3485
rect 6380 3392 6408 3488
rect 9493 3485 9505 3519
rect 9539 3516 9551 3519
rect 9600 3516 9628 3615
rect 9784 3584 9812 3680
rect 10244 3593 10272 3692
rect 10321 3689 10333 3692
rect 10367 3689 10379 3723
rect 10321 3683 10379 3689
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9784 3556 9965 3584
rect 9953 3553 9965 3556
rect 9999 3553 10011 3587
rect 9953 3547 10011 3553
rect 10229 3587 10287 3593
rect 10229 3553 10241 3587
rect 10275 3553 10287 3587
rect 10229 3547 10287 3553
rect 9539 3488 9628 3516
rect 9744 3519 9802 3525
rect 9539 3485 9551 3488
rect 9493 3479 9551 3485
rect 9744 3485 9756 3519
rect 9790 3516 9802 3519
rect 9858 3516 9864 3528
rect 9790 3488 9864 3516
rect 9790 3485 9802 3488
rect 9744 3479 9802 3485
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3485 10563 3519
rect 10505 3479 10563 3485
rect 10520 3448 10548 3479
rect 10152 3420 10548 3448
rect 10152 3392 10180 3420
rect 6362 3340 6368 3392
rect 6420 3340 6426 3392
rect 6457 3383 6515 3389
rect 6457 3349 6469 3383
rect 6503 3380 6515 3383
rect 6546 3380 6552 3392
rect 6503 3352 6552 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 6546 3340 6552 3352
rect 6604 3380 6610 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 6604 3352 9873 3380
rect 6604 3340 6610 3352
rect 9861 3349 9873 3352
rect 9907 3380 9919 3383
rect 10042 3380 10048 3392
rect 9907 3352 10048 3380
rect 9907 3349 9919 3352
rect 9861 3343 9919 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 10134 3340 10140 3392
rect 10192 3340 10198 3392
rect 1104 3290 10856 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 10856 3290
rect 1104 3216 10856 3238
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 4338 3176 4344 3188
rect 3752 3148 4344 3176
rect 3752 3136 3758 3148
rect 4338 3136 4344 3148
rect 4396 3176 4402 3188
rect 5445 3179 5503 3185
rect 4396 3148 4844 3176
rect 4396 3136 4402 3148
rect 3510 3068 3516 3120
rect 3568 3108 3574 3120
rect 4816 3108 4844 3148
rect 5445 3145 5457 3179
rect 5491 3176 5503 3179
rect 10226 3176 10232 3188
rect 5491 3148 10232 3176
rect 5491 3145 5503 3148
rect 5445 3139 5503 3145
rect 5460 3108 5488 3139
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 3568 3080 4016 3108
rect 3568 3068 3574 3080
rect 3528 2981 3556 3068
rect 3602 3000 3608 3052
rect 3660 3000 3666 3052
rect 3694 3000 3700 3052
rect 3752 3000 3758 3052
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2941 3571 2975
rect 3513 2935 3571 2941
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2972 3847 2975
rect 3878 2972 3884 2984
rect 3835 2944 3884 2972
rect 3835 2941 3847 2944
rect 3789 2935 3847 2941
rect 3878 2932 3884 2944
rect 3936 2932 3942 2984
rect 3988 2904 4016 3080
rect 4816 3080 5488 3108
rect 5537 3111 5595 3117
rect 4154 3000 4160 3052
rect 4212 3000 4218 3052
rect 4816 3049 4844 3080
rect 5537 3077 5549 3111
rect 5583 3108 5595 3111
rect 6362 3108 6368 3120
rect 5583 3080 6368 3108
rect 5583 3077 5595 3080
rect 5537 3071 5595 3077
rect 6362 3068 6368 3080
rect 6420 3068 6426 3120
rect 6546 3068 6552 3120
rect 6604 3068 6610 3120
rect 6638 3068 6644 3120
rect 6696 3068 6702 3120
rect 7101 3111 7159 3117
rect 7101 3077 7113 3111
rect 7147 3108 7159 3111
rect 9585 3111 9643 3117
rect 9585 3108 9597 3111
rect 7147 3080 9597 3108
rect 7147 3077 7159 3080
rect 7101 3071 7159 3077
rect 4449 3043 4507 3049
rect 4449 3009 4461 3043
rect 4495 3040 4507 3043
rect 4801 3043 4859 3049
rect 4495 3012 4568 3040
rect 4495 3009 4507 3012
rect 4449 3003 4507 3009
rect 4246 2932 4252 2984
rect 4304 2932 4310 2984
rect 4338 2932 4344 2984
rect 4396 2932 4402 2984
rect 4540 2904 4568 3012
rect 4801 3009 4813 3043
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 7374 3040 7380 3052
rect 5951 3012 7380 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 4614 2932 4620 2984
rect 4672 2932 4678 2984
rect 4890 2932 4896 2984
rect 4948 2932 4954 2984
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2941 5043 2975
rect 4985 2935 5043 2941
rect 5000 2904 5028 2935
rect 5074 2932 5080 2984
rect 5132 2932 5138 2984
rect 5350 2932 5356 2984
rect 5408 2972 5414 2984
rect 7484 2972 7512 3080
rect 9585 3077 9597 3080
rect 9631 3108 9643 3111
rect 10045 3111 10103 3117
rect 10045 3108 10057 3111
rect 9631 3080 10057 3108
rect 9631 3077 9643 3080
rect 9585 3071 9643 3077
rect 10045 3077 10057 3080
rect 10091 3077 10103 3111
rect 10045 3071 10103 3077
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 5408 2944 7512 2972
rect 9508 2972 9536 3003
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 10192 3012 10241 3040
rect 10192 3000 10198 3012
rect 10229 3009 10241 3012
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 9508 2944 9628 2972
rect 5408 2932 5414 2944
rect 9600 2913 9628 2944
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 9950 2972 9956 2984
rect 9732 2944 9956 2972
rect 9732 2932 9738 2944
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 5721 2907 5779 2913
rect 5721 2904 5733 2907
rect 3988 2876 5733 2904
rect 5721 2873 5733 2876
rect 5767 2904 5779 2907
rect 7101 2907 7159 2913
rect 7101 2904 7113 2907
rect 5767 2876 7113 2904
rect 5767 2873 5779 2876
rect 5721 2867 5779 2873
rect 7101 2873 7113 2876
rect 7147 2904 7159 2907
rect 9585 2907 9643 2913
rect 7147 2876 9444 2904
rect 7147 2873 7159 2876
rect 7101 2867 7159 2873
rect 3970 2796 3976 2848
rect 4028 2796 4034 2848
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 4890 2836 4896 2848
rect 4304 2808 4896 2836
rect 4304 2796 4310 2808
rect 4890 2796 4896 2808
rect 4948 2796 4954 2848
rect 5258 2796 5264 2848
rect 5316 2796 5322 2848
rect 6365 2839 6423 2845
rect 6365 2805 6377 2839
rect 6411 2836 6423 2839
rect 6454 2836 6460 2848
rect 6411 2808 6460 2836
rect 6411 2805 6423 2808
rect 6365 2799 6423 2805
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 9306 2796 9312 2848
rect 9364 2796 9370 2848
rect 9416 2836 9444 2876
rect 9585 2873 9597 2907
rect 9631 2873 9643 2907
rect 9585 2867 9643 2873
rect 9861 2907 9919 2913
rect 9861 2873 9873 2907
rect 9907 2904 9919 2907
rect 10226 2904 10232 2916
rect 9907 2876 10232 2904
rect 9907 2873 9919 2876
rect 9861 2867 9919 2873
rect 10226 2864 10232 2876
rect 10284 2864 10290 2916
rect 9769 2839 9827 2845
rect 9769 2836 9781 2839
rect 9416 2808 9781 2836
rect 9769 2805 9781 2808
rect 9815 2805 9827 2839
rect 9769 2799 9827 2805
rect 1104 2746 10856 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 10856 2746
rect 1104 2672 10856 2694
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 4154 2632 4160 2644
rect 3936 2604 4160 2632
rect 3936 2592 3942 2604
rect 4154 2592 4160 2604
rect 4212 2632 4218 2644
rect 5074 2632 5080 2644
rect 4212 2604 5080 2632
rect 4212 2592 4218 2604
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 6454 2632 6460 2644
rect 6196 2604 6460 2632
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 6196 2437 6224 2604
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 6638 2632 6644 2644
rect 6595 2604 6644 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 7374 2592 7380 2644
rect 7432 2592 7438 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 10134 2632 10140 2644
rect 8067 2604 10140 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 8665 2567 8723 2573
rect 8665 2564 8677 2567
rect 6380 2536 8677 2564
rect 6380 2437 6408 2536
rect 8665 2533 8677 2536
rect 8711 2533 8723 2567
rect 8665 2527 8723 2533
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6512 2400 6837 2428
rect 6512 2388 6518 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 8680 2428 8708 2527
rect 9950 2524 9956 2576
rect 10008 2524 10014 2576
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 8680 2400 10149 2428
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3936 2264 4169 2292
rect 3936 2252 3942 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4580 2264 4813 2292
rect 4580 2252 4586 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5224 2264 5457 2292
rect 5224 2252 5230 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 5994 2252 6000 2304
rect 6052 2252 6058 2304
rect 6362 2252 6368 2304
rect 6420 2292 6426 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6420 2264 6653 2292
rect 6420 2252 6426 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 1104 2202 10856 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 10856 2202
rect 1104 2128 10856 2150
<< via1 >>
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 1676 6400 1728 6452
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 3056 6264 3108 6316
rect 10140 6264 10192 6316
rect 2320 6239 2372 6248
rect 2320 6205 2329 6239
rect 2329 6205 2363 6239
rect 2363 6205 2372 6239
rect 2320 6196 2372 6205
rect 2412 6239 2464 6248
rect 2412 6205 2421 6239
rect 2421 6205 2455 6239
rect 2455 6205 2464 6239
rect 2412 6196 2464 6205
rect 9680 6239 9732 6248
rect 9680 6205 9689 6239
rect 9689 6205 9723 6239
rect 9723 6205 9732 6239
rect 9680 6196 9732 6205
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 940 6128 992 6180
rect 2964 6128 3016 6180
rect 9956 6239 10008 6248
rect 9956 6205 9965 6239
rect 9965 6205 9999 6239
rect 9999 6205 10008 6239
rect 9956 6196 10008 6205
rect 10048 6196 10100 6248
rect 10416 6171 10468 6180
rect 10416 6137 10425 6171
rect 10425 6137 10459 6171
rect 10459 6137 10468 6171
rect 10416 6128 10468 6137
rect 9496 6103 9548 6112
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 1676 5899 1728 5908
rect 1676 5865 1685 5899
rect 1685 5865 1719 5899
rect 1719 5865 1728 5899
rect 1676 5856 1728 5865
rect 9496 5856 9548 5908
rect 9864 5856 9916 5908
rect 10232 5899 10284 5908
rect 10232 5865 10241 5899
rect 10241 5865 10275 5899
rect 10275 5865 10284 5899
rect 10232 5856 10284 5865
rect 2320 5788 2372 5840
rect 2780 5788 2832 5840
rect 2964 5788 3016 5840
rect 1768 5652 1820 5704
rect 9680 5720 9732 5772
rect 9772 5720 9824 5772
rect 2320 5584 2372 5636
rect 2780 5627 2832 5636
rect 2780 5593 2789 5627
rect 2789 5593 2823 5627
rect 2823 5593 2832 5627
rect 2780 5584 2832 5593
rect 3516 5584 3568 5636
rect 3056 5516 3108 5568
rect 3148 5516 3200 5568
rect 9312 5559 9364 5568
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 10048 5516 10100 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 848 5312 900 5364
rect 9772 5312 9824 5364
rect 10140 5312 10192 5364
rect 9680 5244 9732 5296
rect 1768 5176 1820 5228
rect 1860 5176 1912 5228
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 9956 5176 10008 5228
rect 9588 5151 9640 5160
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 10232 5108 10284 5160
rect 940 4972 992 5024
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 1860 4768 1912 4820
rect 9496 4768 9548 4820
rect 3148 4700 3200 4752
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 9680 4632 9732 4684
rect 9772 4632 9824 4684
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 2964 4496 3016 4548
rect 10048 4496 10100 4548
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 2228 4471 2280 4480
rect 2228 4437 2237 4471
rect 2237 4437 2271 4471
rect 2271 4437 2280 4471
rect 2228 4428 2280 4437
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 9864 4471 9916 4480
rect 9864 4437 9873 4471
rect 9873 4437 9907 4471
rect 9907 4437 9916 4471
rect 9864 4428 9916 4437
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 1676 4224 1728 4276
rect 2964 4224 3016 4276
rect 3700 4224 3752 4276
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 9772 4224 9824 4276
rect 2228 4156 2280 4208
rect 3056 4156 3108 4208
rect 2320 4088 2372 4140
rect 9956 4088 10008 4140
rect 10048 4131 10100 4140
rect 10048 4097 10057 4131
rect 10057 4097 10091 4131
rect 10091 4097 10100 4131
rect 10048 4088 10100 4097
rect 3516 4020 3568 4072
rect 3884 4020 3936 4072
rect 7380 4020 7432 4072
rect 3148 3995 3200 4004
rect 3148 3961 3157 3995
rect 3157 3961 3191 3995
rect 3191 3961 3200 3995
rect 3148 3952 3200 3961
rect 6644 3952 6696 4004
rect 9864 3952 9916 4004
rect 3608 3884 3660 3936
rect 4252 3884 4304 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 9772 3680 9824 3732
rect 9956 3680 10008 3732
rect 9312 3544 9364 3596
rect 9864 3476 9916 3528
rect 6368 3340 6420 3392
rect 6552 3340 6604 3392
rect 10048 3340 10100 3392
rect 10140 3340 10192 3392
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 3700 3136 3752 3188
rect 4344 3136 4396 3188
rect 3516 3068 3568 3120
rect 10232 3136 10284 3188
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 3884 2932 3936 2984
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 6368 3068 6420 3120
rect 6552 3111 6604 3120
rect 6552 3077 6561 3111
rect 6561 3077 6595 3111
rect 6595 3077 6604 3111
rect 6552 3068 6604 3077
rect 6644 3111 6696 3120
rect 6644 3077 6653 3111
rect 6653 3077 6687 3111
rect 6687 3077 6696 3111
rect 6644 3068 6696 3077
rect 4252 2975 4304 2984
rect 4252 2941 4261 2975
rect 4261 2941 4295 2975
rect 4295 2941 4304 2975
rect 4252 2932 4304 2941
rect 4344 2975 4396 2984
rect 4344 2941 4353 2975
rect 4353 2941 4387 2975
rect 4387 2941 4396 2975
rect 4344 2932 4396 2941
rect 7380 3000 7432 3052
rect 4620 2975 4672 2984
rect 4620 2941 4629 2975
rect 4629 2941 4663 2975
rect 4663 2941 4672 2975
rect 4620 2932 4672 2941
rect 4896 2975 4948 2984
rect 4896 2941 4905 2975
rect 4905 2941 4939 2975
rect 4939 2941 4948 2975
rect 4896 2932 4948 2941
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 5356 2932 5408 2984
rect 10140 3000 10192 3052
rect 9680 2932 9732 2984
rect 9956 2975 10008 2984
rect 9956 2941 9965 2975
rect 9965 2941 9999 2975
rect 9999 2941 10008 2975
rect 9956 2932 10008 2941
rect 3976 2839 4028 2848
rect 3976 2805 3985 2839
rect 3985 2805 4019 2839
rect 4019 2805 4028 2839
rect 3976 2796 4028 2805
rect 4252 2796 4304 2848
rect 4896 2796 4948 2848
rect 5264 2839 5316 2848
rect 5264 2805 5273 2839
rect 5273 2805 5307 2839
rect 5307 2805 5316 2839
rect 5264 2796 5316 2805
rect 6460 2796 6512 2848
rect 9312 2839 9364 2848
rect 9312 2805 9321 2839
rect 9321 2805 9355 2839
rect 9355 2805 9364 2839
rect 9312 2796 9364 2805
rect 10232 2864 10284 2916
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 3884 2592 3936 2644
rect 4160 2592 4212 2644
rect 5080 2592 5132 2644
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 6460 2592 6512 2644
rect 6644 2592 6696 2644
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 10140 2592 10192 2644
rect 6460 2388 6512 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 9956 2567 10008 2576
rect 9956 2533 9965 2567
rect 9965 2533 9999 2567
rect 9999 2533 10008 2567
rect 9956 2524 10008 2533
rect 3884 2252 3936 2304
rect 4528 2252 4580 2304
rect 5172 2252 5224 2304
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 6368 2252 6420 2304
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
<< metal2 >>
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6905 1532 7142
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1688 6458 1716 7346
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 938 6216 994 6225
rect 938 6151 940 6160
rect 992 6151 994 6160
rect 940 6122 992 6128
rect 1688 5914 1716 6258
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 2332 5846 2360 6190
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 846 5400 902 5409
rect 846 5335 848 5344
rect 900 5335 902 5344
rect 848 5306 900 5312
rect 1780 5234 1808 5646
rect 2320 5636 2372 5642
rect 2424 5624 2452 6190
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2976 5846 3004 6122
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2792 5642 2820 5782
rect 2372 5596 2452 5624
rect 2780 5636 2832 5642
rect 2320 5578 2372 5584
rect 2780 5578 2832 5584
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4865 980 4966
rect 938 4856 994 4865
rect 1872 4826 1900 5170
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 938 4791 994 4800
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4185 1532 4422
rect 1688 4282 1716 4558
rect 2332 4486 2360 5578
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2976 4554 3004 5782
rect 3068 5574 3096 6258
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9772 6248 9824 6254
rect 9956 6248 10008 6254
rect 9772 6190 9824 6196
rect 9876 6208 9956 6236
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 9508 5914 9536 6054
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9692 5778 9720 6190
rect 9784 5778 9812 6190
rect 9876 5914 9904 6208
rect 9956 6190 10008 6196
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 2240 4214 2268 4422
rect 2228 4208 2280 4214
rect 1490 4176 1546 4185
rect 2228 4150 2280 4156
rect 2332 4146 2360 4422
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2976 4282 3004 4490
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 3068 4214 3096 5510
rect 3160 4758 3188 5510
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 1490 4111 1546 4120
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 3160 4010 3188 4694
rect 3528 4078 3556 5578
rect 9312 5568 9364 5574
rect 9310 5536 9312 5545
rect 9364 5536 9366 5545
rect 7610 5468 7918 5477
rect 9310 5471 9366 5480
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 9692 5302 9720 5714
rect 9784 5370 9812 5714
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 9324 4865 9352 4966
rect 9310 4856 9366 4865
rect 9508 4826 9536 5170
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9310 4791 9366 4800
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 3528 3126 3556 4014
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3620 3058 3648 3878
rect 3712 3194 3740 4218
rect 9324 4185 9352 4422
rect 9310 4176 9366 4185
rect 9310 4111 9366 4120
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3712 3058 3740 3130
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3896 2990 3924 4014
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 3896 2650 3924 2926
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3988 2446 4016 2790
rect 4172 2650 4200 2994
rect 4264 2990 4292 3878
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4356 2990 4384 3130
rect 6380 3126 6408 3334
rect 6564 3126 6592 3334
rect 6656 3126 6684 3946
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4896 2984 4948 2990
rect 5080 2984 5132 2990
rect 4986 2952 5042 2961
rect 4948 2932 4986 2938
rect 4896 2926 4986 2932
rect 4264 2854 4292 2926
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4632 2446 4660 2926
rect 4908 2910 4986 2926
rect 4908 2854 4936 2910
rect 5356 2984 5408 2990
rect 5132 2944 5356 2972
rect 5080 2926 5132 2932
rect 5356 2926 5408 2932
rect 4986 2887 5042 2896
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 5092 2650 5120 2926
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5276 2446 5304 2790
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6380 2310 6408 3062
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6472 2650 6500 2790
rect 6656 2650 6684 3062
rect 7392 3058 7420 4014
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9324 3505 9352 3538
rect 9310 3496 9366 3505
rect 9310 3431 9366 3440
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 7392 2650 7420 2994
rect 9600 2972 9628 5102
rect 9784 4690 9812 5306
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9692 4282 9720 4626
rect 9784 4282 9812 4626
rect 9876 4486 9904 5850
rect 10060 5574 10088 6190
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9968 4622 9996 5170
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9784 3738 9812 4218
rect 9876 4010 9904 4422
rect 9968 4146 9996 4558
rect 10060 4554 10088 5510
rect 10152 5370 10180 6258
rect 10244 5914 10272 7346
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10428 6905 10456 7142
rect 10414 6896 10470 6905
rect 10414 6831 10470 6840
rect 10414 6216 10470 6225
rect 10414 6151 10416 6160
rect 10468 6151 10470 6160
rect 10416 6122 10468 6128
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 10060 4146 10088 4490
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9876 3534 9904 3946
rect 9968 3738 9996 4082
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10060 3398 10088 4082
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 3058 10180 3334
rect 10244 3194 10272 5102
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 9680 2984 9732 2990
rect 9600 2961 9680 2972
rect 9586 2952 9680 2961
rect 9642 2944 9680 2952
rect 9680 2926 9732 2932
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9586 2887 9642 2896
rect 9312 2848 9364 2854
rect 9310 2816 9312 2825
rect 9364 2816 9366 2825
rect 9310 2751 9366 2760
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 9968 2582 9996 2926
rect 10152 2650 10180 2994
rect 10244 2922 10272 3130
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 6460 2440 6512 2446
rect 7196 2440 7248 2446
rect 6460 2382 6512 2388
rect 7116 2400 7196 2428
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 3896 800 3924 2246
rect 4540 800 4568 2246
rect 5184 800 5212 2246
rect 6012 1170 6040 2246
rect 5828 1142 6040 1170
rect 5828 800 5856 1142
rect 6472 800 6500 2382
rect 7116 800 7144 2400
rect 7196 2382 7248 2388
rect 7840 2440 7892 2446
rect 8484 2440 8536 2446
rect 7892 2400 8064 2428
rect 7840 2382 7892 2388
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 7760 870 7880 898
rect 7760 800 7788 870
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 7852 762 7880 870
rect 8036 762 8064 2400
rect 8404 2400 8484 2428
rect 8404 800 8432 2400
rect 8484 2382 8536 2388
rect 7852 734 8064 762
rect 8390 0 8446 800
<< via2 >>
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 1490 6840 1546 6896
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 938 6180 994 6216
rect 938 6160 940 6180
rect 940 6160 992 6180
rect 992 6160 994 6180
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 846 5364 902 5400
rect 846 5344 848 5364
rect 848 5344 900 5364
rect 900 5344 902 5364
rect 938 4800 994 4856
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 1490 4120 1546 4176
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 9310 5516 9312 5536
rect 9312 5516 9364 5536
rect 9364 5516 9366 5536
rect 9310 5480 9366 5516
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 9310 4800 9366 4856
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 9310 4120 9366 4176
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 4986 2896 5042 2952
rect 9310 3440 9366 3496
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 10414 6840 10470 6896
rect 10414 6180 10470 6216
rect 10414 6160 10416 6180
rect 10416 6160 10468 6180
rect 10468 6160 10470 6180
rect 9586 2896 9642 2952
rect 9310 2796 9312 2816
rect 9312 2796 9364 2816
rect 9364 2796 9366 2816
rect 9310 2760 9366 2796
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
<< metal3 >>
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 10409 6898 10475 6901
rect 11200 6898 12000 6928
rect 10409 6896 12000 6898
rect 10409 6840 10414 6896
rect 10470 6840 12000 6896
rect 10409 6838 12000 6840
rect 10409 6835 10475 6838
rect 11200 6808 12000 6838
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 0 6218 800 6248
rect 933 6218 999 6221
rect 0 6216 999 6218
rect 0 6160 938 6216
rect 994 6160 999 6216
rect 0 6158 999 6160
rect 0 6128 800 6158
rect 933 6155 999 6158
rect 10409 6218 10475 6221
rect 11200 6218 12000 6248
rect 10409 6216 12000 6218
rect 10409 6160 10414 6216
rect 10470 6160 12000 6216
rect 10409 6158 12000 6160
rect 10409 6155 10475 6158
rect 11200 6128 12000 6158
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 0 5538 800 5568
rect 9305 5538 9371 5541
rect 11200 5538 12000 5568
rect 0 5448 858 5538
rect 9305 5536 12000 5538
rect 9305 5480 9310 5536
rect 9366 5480 12000 5536
rect 9305 5478 12000 5480
rect 9305 5475 9371 5478
rect 798 5405 858 5448
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 11200 5448 12000 5478
rect 7606 5407 7922 5408
rect 798 5400 907 5405
rect 798 5344 846 5400
rect 902 5344 907 5400
rect 798 5342 907 5344
rect 841 5339 907 5342
rect 1946 4928 2262 4929
rect 0 4858 800 4888
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 9305 4858 9371 4861
rect 11200 4858 12000 4888
rect 9305 4856 12000 4858
rect 9305 4800 9310 4856
rect 9366 4800 12000 4856
rect 9305 4798 12000 4800
rect 9305 4795 9371 4798
rect 11200 4768 12000 4798
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 0 4178 800 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 904 4118
rect 1485 4115 1551 4118
rect 9305 4178 9371 4181
rect 11200 4178 12000 4208
rect 9305 4176 12000 4178
rect 9305 4120 9310 4176
rect 9366 4120 12000 4176
rect 9305 4118 12000 4120
rect 9305 4115 9371 4118
rect 11200 4088 12000 4118
rect 798 4084 904 4088
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 9305 3498 9371 3501
rect 11200 3498 12000 3528
rect 9305 3496 12000 3498
rect 9305 3440 9310 3496
rect 9366 3440 12000 3496
rect 9305 3438 12000 3440
rect 9305 3435 9371 3438
rect 11200 3408 12000 3438
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 4981 2954 5047 2957
rect 9581 2954 9647 2957
rect 4981 2952 9647 2954
rect 4981 2896 4986 2952
rect 5042 2896 9586 2952
rect 9642 2896 9647 2952
rect 4981 2894 9647 2896
rect 4981 2891 5047 2894
rect 9581 2891 9647 2894
rect 9305 2818 9371 2821
rect 11200 2818 12000 2848
rect 9305 2816 12000 2818
rect 9305 2760 9310 2816
rect 9366 2760 12000 2816
rect 9305 2758 12000 2760
rect 9305 2755 9371 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 11200 2728 12000 2758
rect 6946 2687 7262 2688
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
<< via3 >>
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
<< metal4 >>
rect 1944 9280 2264 9840
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 9824 2924 9840
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 9280 7264 9840
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 9824 7924 9840
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7604 7648 7924 8672
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
<< via4 >>
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1986 3058 2222 3294
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 2646 3718 2882 3954
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 6986 3058 7222 3294
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 7646 3718 7882 3954
<< metal5 >>
rect 1056 8954 10904 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 10904 8954
rect 1056 8676 10904 8718
rect 1056 8294 10904 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 10904 8294
rect 1056 8016 10904 8058
rect 1056 3954 10904 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 10904 3954
rect 1056 3676 10904 3718
rect 1056 3294 10904 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 10904 3294
rect 1056 3016 10904 3058
use sky130_fd_sc_hd__nor4_1  _00_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 9568 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  _01_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 5336 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _02_
timestamp 1707688321
transform -1 0 4048 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _03_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 3312 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _04_
timestamp 1707688321
transform -1 0 4692 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _05_
timestamp 1707688321
transform -1 0 2576 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _06_
timestamp 1707688321
transform -1 0 2944 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _07_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 9568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _08_
timestamp 1707688321
transform 1 0 9476 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _09_
timestamp 1707688321
transform -1 0 7268 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _10_
timestamp 1707688321
transform -1 0 3036 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _11_
timestamp 1707688321
transform -1 0 10304 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _12_
timestamp 1707688321
transform -1 0 3496 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _13_
timestamp 1707688321
transform -1 0 10304 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _14_
timestamp 1707688321
transform 1 0 9568 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 10304 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  fanout21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 1707688321
transform -1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout24
timestamp 1707688321
transform -1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1707688321
transform -1 0 6072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout26
timestamp 1707688321
transform -1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1707688321
transform -1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout28
timestamp 1707688321
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1707688321
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_42
timestamp 1707688321
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_49
timestamp 1707688321
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_63
timestamp 1707688321
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_76
timestamp 1707688321
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1707688321
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_93
timestamp 1707688321
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_100
timestamp 1707688321
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1707688321
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_15
timestamp 1707688321
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_23
timestamp 1707688321
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1707688321
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_67
timestamp 1707688321
transform 1 0 7268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_79
timestamp 1707688321
transform 1 0 8372 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_87
timestamp 1707688321
transform 1 0 9108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_101
timestamp 1707688321
transform 1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1707688321
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1707688321
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1707688321
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1707688321
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1707688321
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_53
timestamp 1707688321
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_59
timestamp 1707688321
transform 1 0 6532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_71
timestamp 1707688321
transform 1 0 7636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1707688321
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_85
timestamp 1707688321
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1707688321
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_11
timestamp 1707688321
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_24
timestamp 1707688321
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_36
timestamp 1707688321
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_48
timestamp 1707688321
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1707688321
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1707688321
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1707688321
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_7
timestamp 1707688321
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_20
timestamp 1707688321
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1707688321
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1707688321
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1707688321
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1707688321
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1707688321
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 1707688321
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_100
timestamp 1707688321
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_11
timestamp 1707688321
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_23
timestamp 1707688321
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_35
timestamp 1707688321
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_47
timestamp 1707688321
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1707688321
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1707688321
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1707688321
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_81
timestamp 1707688321
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_87
timestamp 1707688321
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_100
timestamp 1707688321
transform 1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 1707688321
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1707688321
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1707688321
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1707688321
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1707688321
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1707688321
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1707688321
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1707688321
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_85
timestamp 1707688321
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_100
timestamp 1707688321
transform 1 0 10304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_7
timestamp 1707688321
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_21
timestamp 1707688321
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_33
timestamp 1707688321
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_45
timestamp 1707688321
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1707688321
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1707688321
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1707688321
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_81
timestamp 1707688321
transform 1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_89
timestamp 1707688321
transform 1 0 9292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_98
timestamp 1707688321
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1707688321
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1707688321
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1707688321
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1707688321
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1707688321
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1707688321
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1707688321
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1707688321
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1707688321
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1707688321
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_97
timestamp 1707688321
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_7
timestamp 1707688321
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_19
timestamp 1707688321
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_31
timestamp 1707688321
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_43
timestamp 1707688321
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1707688321
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1707688321
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1707688321
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1707688321
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_93
timestamp 1707688321
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1707688321
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1707688321
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1707688321
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1707688321
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1707688321
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1707688321
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1707688321
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1707688321
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1707688321
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1707688321
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_97
timestamp 1707688321
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1707688321
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1707688321
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1707688321
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1707688321
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1707688321
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1707688321
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1707688321
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1707688321
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1707688321
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_93
timestamp 1707688321
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_101
timestamp 1707688321
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1707688321
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1707688321
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1707688321
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1707688321
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1707688321
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1707688321
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1707688321
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1707688321
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1707688321
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1707688321
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_97
timestamp 1707688321
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1707688321
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1707688321
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1707688321
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_29
timestamp 1707688321
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 1707688321
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1707688321
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1707688321
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1707688321
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_81
timestamp 1707688321
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_85
timestamp 1707688321
transform 1 0 8924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_97
timestamp 1707688321
transform 1 0 10028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1707688321
transform -1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1707688321
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1707688321
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1707688321
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1707688321
transform -1 0 9568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1707688321
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1707688321
transform -1 0 9568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1707688321
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1707688321
transform -1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1707688321
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1707688321
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1707688321
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1707688321
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1707688321
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1707688321
transform -1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1707688321
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1707688321
transform -1 0 9568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1707688321
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_14
timestamp 1707688321
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1707688321
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_15
timestamp 1707688321
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1707688321
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_16
timestamp 1707688321
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1707688321
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_17
timestamp 1707688321
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1707688321
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_18
timestamp 1707688321
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1707688321
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_19
timestamp 1707688321
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1707688321
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_20
timestamp 1707688321
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1707688321
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_21
timestamp 1707688321
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1707688321
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_22
timestamp 1707688321
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1707688321
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_23
timestamp 1707688321
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1707688321
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_24
timestamp 1707688321
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1707688321
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_25
timestamp 1707688321
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1707688321
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_26
timestamp 1707688321
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1707688321
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_27
timestamp 1707688321
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1707688321
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp 1707688321
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp 1707688321
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_31
timestamp 1707688321
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_32
timestamp 1707688321
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_33
timestamp 1707688321
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_34
timestamp 1707688321
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_35
timestamp 1707688321
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_36
timestamp 1707688321
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_37
timestamp 1707688321
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_38
timestamp 1707688321
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_39
timestamp 1707688321
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_40
timestamp 1707688321
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_41
timestamp 1707688321
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_42
timestamp 1707688321
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_43
timestamp 1707688321
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_44
timestamp 1707688321
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_45
timestamp 1707688321
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_46
timestamp 1707688321
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_47
timestamp 1707688321
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_48
timestamp 1707688321
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_49
timestamp 1707688321
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_50
timestamp 1707688321
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_51
timestamp 1707688321
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal4 s 2604 2128 2924 9840 0 FreeSans 1920 90 0 0 VGND
port 18 nsew ground bidirectional
flabel metal4 s 7604 2128 7924 9840 0 FreeSans 1920 90 0 0 VGND
port 18 nsew ground bidirectional
flabel metal5 s 1056 3676 10904 3996 0 FreeSans 2560 0 0 0 VGND
port 18 nsew ground bidirectional
flabel metal5 s 1056 8676 10904 8996 0 FreeSans 2560 0 0 0 VGND
port 18 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6944 2128 7264 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3016 10904 3336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8016 10904 8336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 otrip[0]
port 22 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 otrip[1]
port 21 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 otrip[2]
port 20 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 otrip[3]
port 19 nsew signal input
flabel metal3 s 11200 2728 12000 2848 0 FreeSans 480 0 0 0 otrip_decoded[0]
port 17 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 otrip_decoded[10]
port 7 nsew signal output
flabel metal3 s 11200 3408 12000 3528 0 FreeSans 480 0 0 0 otrip_decoded[11]
port 6 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 otrip_decoded[12]
port 5 nsew signal output
flabel metal3 s 11200 4768 12000 4888 0 FreeSans 480 0 0 0 otrip_decoded[13]
port 4 nsew signal output
flabel metal3 s 11200 6808 12000 6928 0 FreeSans 480 0 0 0 otrip_decoded[14]
port 3 nsew signal output
flabel metal3 s 11200 4088 12000 4208 0 FreeSans 480 0 0 0 otrip_decoded[15]
port 2 nsew signal output
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 otrip_decoded[1]
port 16 nsew signal output
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 otrip_decoded[2]
port 15 nsew signal output
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 otrip_decoded[3]
port 14 nsew signal output
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 otrip_decoded[4]
port 13 nsew signal output
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 otrip_decoded[5]
port 12 nsew signal output
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 otrip_decoded[6]
port 11 nsew signal output
flabel metal3 s 11200 6128 12000 6248 0 FreeSans 480 0 0 0 otrip_decoded[7]
port 10 nsew signal output
flabel metal3 s 11200 5448 12000 5568 0 FreeSans 480 0 0 0 otrip_decoded[8]
port 9 nsew signal output
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 otrip_decoded[9]
port 8 nsew signal output
rlabel metal1 5980 9792 5980 9792 0 VGND
rlabel metal1 5980 9248 5980 9248 0 VPWR
rlabel metal1 6532 2278 6532 2278 0 net1
rlabel metal2 10258 6630 10258 6630 0 net10
rlabel metal2 9706 4454 9706 4454 0 net11
rlabel metal2 5290 2618 5290 2618 0 net12
rlabel metal2 4002 2618 4002 2618 0 net13
rlabel metal1 2070 4250 2070 4250 0 net14
rlabel metal2 4646 2686 4646 2686 0 net15
rlabel metal2 1702 6086 1702 6086 0 net16
rlabel metal1 1978 4794 1978 4794 0 net17
rlabel metal1 10212 5338 10212 5338 0 net18
rlabel metal1 9522 5780 9522 5780 0 net19
rlabel metal1 8970 4046 8970 4046 0 net2
rlabel metal1 6210 2516 6210 2516 0 net20
rlabel metal1 9844 2958 9844 2958 0 net21
rlabel metal1 6624 2618 6624 2618 0 net22
rlabel metal1 8372 3094 8372 3094 0 net23
rlabel metal1 9844 5678 9844 5678 0 net24
rlabel metal1 8280 2890 8280 2890 0 net25
rlabel metal1 9844 5746 9844 5746 0 net26
rlabel metal1 10074 5134 10074 5134 0 net27
rlabel metal1 6532 3366 6532 3366 0 net28
rlabel metal1 9108 2618 9108 2618 0 net3
rlabel metal1 6394 2482 6394 2482 0 net4
rlabel metal1 9522 2992 9522 2992 0 net5
rlabel metal1 1932 6426 1932 6426 0 net6
rlabel metal1 9568 3502 9568 3502 0 net7
rlabel metal1 1748 5202 1748 5202 0 net8
rlabel metal1 9568 4794 9568 4794 0 net9
rlabel metal2 6486 1588 6486 1588 0 otrip[0]
rlabel metal2 7130 1588 7130 1588 0 otrip[1]
rlabel metal2 7774 823 7774 823 0 otrip[2]
rlabel metal2 8418 1588 8418 1588 0 otrip[3]
rlabel via2 9338 2805 9338 2805 0 otrip_decoded[0]
rlabel metal3 1096 6868 1096 6868 0 otrip_decoded[10]
rlabel metal1 9338 3638 9338 3638 0 otrip_decoded[11]
rlabel metal1 1196 5338 1196 5338 0 otrip_decoded[12]
rlabel metal2 9338 4913 9338 4913 0 otrip_decoded[13]
rlabel metal2 10442 7021 10442 7021 0 otrip_decoded[14]
rlabel metal2 9338 4301 9338 4301 0 otrip_decoded[15]
rlabel metal2 5198 1520 5198 1520 0 otrip_decoded[1]
rlabel metal2 3910 1520 3910 1520 0 otrip_decoded[2]
rlabel metal3 751 4148 751 4148 0 otrip_decoded[3]
rlabel metal2 4554 1520 4554 1520 0 otrip_decoded[4]
rlabel metal3 820 6188 820 6188 0 otrip_decoded[5]
rlabel metal3 820 4828 820 4828 0 otrip_decoded[6]
rlabel via2 10442 6171 10442 6171 0 otrip_decoded[7]
rlabel via2 9338 5525 9338 5525 0 otrip_decoded[8]
rlabel metal2 5842 959 5842 959 0 otrip_decoded[9]
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
