** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/sky130_ajc_ip__overvoltage.sch
.subckt sky130_ajc_ip__overvoltage avdd avss dvdd dvss vbg_1v2 ovout itest otrip[3] otrip[2] otrip[1] otrip[0] vin ena isrc_sel
+ ibg_200n
*.PININFO avdd:I avss:I dvdd:I dvss:I vbg_1v2:I otrip[3:0]:I ena:I isrc_sel:I ibg_200n:I vin:O ovout:O itest:O
xIana otrip_decoded_15_ otrip_decoded_14_ otrip_decoded_13_ otrip_decoded_12_ otrip_decoded_11_ otrip_decoded_10_ otrip_decoded_9_
+ otrip_decoded_8_ otrip_decoded_7_ otrip_decoded_6_ otrip_decoded_5_ otrip_decoded_4_ otrip_decoded_3_ otrip_decoded_2_ otrip_decoded_1_
+ otrip_decoded_0_ vbg_1v2 ena avdd avss dvdd isrc_sel dvss vin itest ibg_200n ovout overvoltage_ana
**** begin user architecture code



*XSPICE CO-SIM netlist
.include overvoltage_dig.out.spice

r0 otrip[0] otrip0 1
r1 otrip[1] otrip1 1
r2 otrip[2] otrip2 1
r3 otrip[3] otrip3 1

xiovervoltage_dig dvss dvdd
+otrip0 otrip1 otrip2 otrip3
+otrip_decoded_0_
+otrip_decoded_10_ otrip_decoded_11_ otrip_decoded_12_ otrip_decoded_13_ otrip_decoded_14_ otrip_decoded_15_
+otrip_decoded_1_ otrip_decoded_2_ otrip_decoded_3_ otrip_decoded_4_ otrip_decoded_5_ otrip_decoded_6_ otrip_decoded_7_
+otrip_decoded_8_ otrip_decoded_9_
+overvoltage_dig



**** end user architecture code
.ends

* expanding   symbol:  xschem/overvoltage_ana.sym # of pins=12
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/overvoltage_ana.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/overvoltage_ana.sch
.subckt overvoltage_ana otrip_decoded[15] otrip_decoded[14] otrip_decoded[13] otrip_decoded[12] otrip_decoded[11]
+ otrip_decoded[10] otrip_decoded[9] otrip_decoded[8] otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[4] otrip_decoded[3]
+ otrip_decoded[2] otrip_decoded[1] otrip_decoded[0] vbg_1v2 ena avdd avss dvdd isrc_sel dvss vin itest ibg_200n ovout
*.PININFO vbg_1v2:I avdd:I avss:I dvdd:I dvss:I ena:I isrc_sel:I ibg_200n:I ovout:O itest:O otrip_decoded[15:0]:I vin:O
XR1 dcomp_filt dcomp avss sky130_fd_pr__res_xhigh_po W=2 L=1000 mult=1 m=1
xIlvls4 dcomp_filt dvdd avss avss avdd avdd net2 sky130_fd_sc_hvl__lsbufhv2lv_1
XC1 dcomp_filt avss sky130_fd_pr__cap_mim_m3_1 W=30 L=30 m=3
XC2 dcomp_filt avss sky130_fd_pr__cap_mim_m3_2 W=30 L=30 m=3
xIlvls0[15] otrip_decoded[15] dvdd avss avss avdd avdd otrip_decoded_avdd[15] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[14] otrip_decoded[14] dvdd avss avss avdd avdd otrip_decoded_avdd[14] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[13] otrip_decoded[13] dvdd avss avss avdd avdd otrip_decoded_avdd[13] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[12] otrip_decoded[12] dvdd avss avss avdd avdd otrip_decoded_avdd[12] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[11] otrip_decoded[11] dvdd avss avss avdd avdd otrip_decoded_avdd[11] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[10] otrip_decoded[10] dvdd avss avss avdd avdd otrip_decoded_avdd[10] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[9] otrip_decoded[9] dvdd avss avss avdd avdd otrip_decoded_avdd[9] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[8] otrip_decoded[8] dvdd avss avss avdd avdd otrip_decoded_avdd[8] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[7] otrip_decoded[7] dvdd avss avss avdd avdd otrip_decoded_avdd[7] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[6] otrip_decoded[6] dvdd avss avss avdd avdd otrip_decoded_avdd[6] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[5] otrip_decoded[5] dvdd avss avss avdd avdd otrip_decoded_avdd[5] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[4] otrip_decoded[4] dvdd avss avss avdd avdd otrip_decoded_avdd[4] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[3] otrip_decoded[3] dvdd avss avss avdd avdd otrip_decoded_avdd[3] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[2] otrip_decoded[2] dvdd avss avss avdd avdd otrip_decoded_avdd[2] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[1] otrip_decoded[1] dvdd avss avss avdd avdd otrip_decoded_avdd[1] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[0] otrip_decoded[0] dvdd avss avss avdd avdd otrip_decoded_avdd[0] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls1 ena dvdd avss avss avdd avdd ena_avdd sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls2 isrc_sel dvdd avss avss avdd avdd isrc_sel_avdd sky130_fd_sc_hvl__lsbuflv2hv_1
xIrsmux avdd vin otrip_decoded_avdd[15] otrip_decoded_avdd[14] otrip_decoded_avdd[13] otrip_decoded_avdd[12]
+ otrip_decoded_avdd[11] otrip_decoded_avdd[10] otrip_decoded_avdd[9] otrip_decoded_avdd[8] otrip_decoded_avdd[7] otrip_decoded_avdd[6]
+ otrip_decoded_avdd[5] otrip_decoded_avdd[4] otrip_decoded_avdd[3] otrip_decoded_avdd[2] otrip_decoded_avdd[1] otrip_decoded_avdd[0] dvdd dvss ena_avdd
+ avss rstring_mux
xIcomp avdd ibias dcomp ena_avdd vbg_1v2 vin avss comparator
xIbiasgen avdd itest ibias ibg_200n vbg_1v2 isrc_sel_avdd ena_avdd avss ibias_gen
xIinv3 net2 dvss dvss dvdd dvdd net1 sky130_fd_sc_hd__inv_4
xIinv4 net1 dvss dvss dvdd dvdd ovout sky130_fd_sc_hd__inv_16
.ends


* expanding   symbol:  rstring_mux.sym # of pins=7
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/rstring_mux.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/rstring_mux.sch
.subckt rstring_mux avdd vout otrip_decoded_avdd[15] otrip_decoded_avdd[14] otrip_decoded_avdd[13] otrip_decoded_avdd[12]
+ otrip_decoded_avdd[11] otrip_decoded_avdd[10] otrip_decoded_avdd[9] otrip_decoded_avdd[8] otrip_decoded_avdd[7] otrip_decoded_avdd[6]
+ otrip_decoded_avdd[5] otrip_decoded_avdd[4] otrip_decoded_avdd[3] otrip_decoded_avdd[2] otrip_decoded_avdd[1] otrip_decoded_avdd[0] dvdd dvss ena avss
*.PININFO avdd:I avss:I vout:O ena:I otrip_decoded_avdd[15:0]:I dvss:I dvdd:I
XR1 net3 net4 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR2 net4 net5 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR0 net1 net3 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR3 net5 net6 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR4 net6 net7 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR5 net7 net8 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR6 net8 net9 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR7 net9 net10 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR8 net10 net11 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR9 net11 net12 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR10 net12 net13 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR11 net13 net14 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR12 net14 net15 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR13 net15 net16 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR14 net16 net17 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR15 net17 net18 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR16 net18 net19 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR17 net19 net20 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR18 net20 net21 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR19 net21 net22 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR20 net22 net23 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR21 net23 net24 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR22 net24 vtrip15 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR23 vtrip15 vtrip14 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR24 vtrip14 vtrip13 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR25 vtrip13 vtrip12 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR26 vtrip12 vtrip11 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR27 vtrip11 vtrip10 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR28 vtrip10 vtrip9 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR29 vtrip9 vtrip8 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR30 vtrip8 vtrip7 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR31 vtrip7 vtrip6 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR32 vtrip6 vtrip5 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR33 vtrip5 vtrip4 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR34 vtrip4 vtrip3 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR35 vtrip3 vtrip2 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR36 vtrip2 vtrip1 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR37 vtrip1 vtrip0 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR38 vtrip0 net25 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR39 net25 net26 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR40 net26 net27 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR41 net27 net28 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR42 net28 net29 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR43 net29 net30 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR44 net30 net31 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR45 net31 net32 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR46 net32 net33 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR47 net33 net34 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR48 net34 net35 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR49 net35 net36 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR50 net36 net37 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR51 net37 net38 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR52 net38 net39 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR53 net39 net40 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR54 net40 net41 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR55 net41 net42 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR56 net42 net43 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR57 net43 net44 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR58 net44 net45 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR59 net45 net46 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR60 net46 net47 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR61 net47 net48 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR62 net48 net49 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR63 net49 net50 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR64 net50 net51 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR65 net51 net52 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR66 net52 net53 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR67 net53 net54 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR68 net54 net55 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR69 net55 net56 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XMtp[15] vtrip15 otrip_decoded_b_avdd[15] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[14] vtrip14 otrip_decoded_b_avdd[14] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[13] vtrip13 otrip_decoded_b_avdd[13] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[12] vtrip12 otrip_decoded_b_avdd[12] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[11] vtrip11 otrip_decoded_b_avdd[11] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[10] vtrip10 otrip_decoded_b_avdd[10] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[9] vtrip9 otrip_decoded_b_avdd[9] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[8] vtrip8 otrip_decoded_b_avdd[8] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[7] vtrip7 otrip_decoded_b_avdd[7] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[6] vtrip6 otrip_decoded_b_avdd[6] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[5] vtrip5 otrip_decoded_b_avdd[5] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[4] vtrip4 otrip_decoded_b_avdd[4] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[3] vtrip3 otrip_decoded_b_avdd[3] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[2] vtrip2 otrip_decoded_b_avdd[2] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[1] vtrip1 otrip_decoded_b_avdd[1] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[0] vtrip0 otrip_decoded_b_avdd[0] vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[15] vout otrip_decoded_avdd[15] vtrip15 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[14] vout otrip_decoded_avdd[14] vtrip14 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[13] vout otrip_decoded_avdd[13] vtrip13 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[12] vout otrip_decoded_avdd[12] vtrip12 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[11] vout otrip_decoded_avdd[11] vtrip11 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[10] vout otrip_decoded_avdd[10] vtrip10 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[9] vout otrip_decoded_avdd[9] vtrip9 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[8] vout otrip_decoded_avdd[8] vtrip8 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[7] vout otrip_decoded_avdd[7] vtrip7 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[6] vout otrip_decoded_avdd[6] vtrip6 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[5] vout otrip_decoded_avdd[5] vtrip5 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[4] vout otrip_decoded_avdd[4] vtrip4 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[3] vout otrip_decoded_avdd[3] vtrip3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[2] vout otrip_decoded_avdd[2] vtrip2 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[1] vout otrip_decoded_avdd[1] vtrip1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[0] vout otrip_decoded_avdd[0] vtrip0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMena net1 ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=16
XR70 net56 net2 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR71 net2 net57 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR72 net57 net58 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR73 net58 net59 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR74 net59 net60 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR75 net60 net61 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR76 net61 net62 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR77 net62 net63 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR78 net63 net64 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR79 net64 net65 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR80 net65 net66 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR81 net66 net67 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR82 net67 net68 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR83 net68 net69 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR84 net69 net70 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR85 net70 net71 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR86 net71 net72 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR87 net72 net73 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR88 net73 net74 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR89 net74 net75 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR90 net75 net76 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR91 net76 net77 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR92 net77 net78 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR93 net78 net79 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR94 net79 net80 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR95 net80 net81 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR96 net81 net82 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR97 net82 net83 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR98 net83 net84 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR99 net84 net85 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR100 net85 net86 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR101 net86 net87 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR102 net87 net88 avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
XR103 net88 avdd avss sky130_fd_pr__res_xhigh_po W=2 L=25 mult=1 m=1
xIinv[15] otrip_decoded_avdd[15] VGND VNB VPB VPWR otrip_decoded_b_avdd[15] sky130_fd_sc_hvl__inv_1
xIinv[14] otrip_decoded_avdd[14] VGND VNB VPB VPWR otrip_decoded_b_avdd[14] sky130_fd_sc_hvl__inv_1
xIinv[13] otrip_decoded_avdd[13] VGND VNB VPB VPWR otrip_decoded_b_avdd[13] sky130_fd_sc_hvl__inv_1
xIinv[12] otrip_decoded_avdd[12] VGND VNB VPB VPWR otrip_decoded_b_avdd[12] sky130_fd_sc_hvl__inv_1
xIinv[11] otrip_decoded_avdd[11] VGND VNB VPB VPWR otrip_decoded_b_avdd[11] sky130_fd_sc_hvl__inv_1
xIinv[10] otrip_decoded_avdd[10] VGND VNB VPB VPWR otrip_decoded_b_avdd[10] sky130_fd_sc_hvl__inv_1
xIinv[9] otrip_decoded_avdd[9] VGND VNB VPB VPWR otrip_decoded_b_avdd[9] sky130_fd_sc_hvl__inv_1
xIinv[8] otrip_decoded_avdd[8] VGND VNB VPB VPWR otrip_decoded_b_avdd[8] sky130_fd_sc_hvl__inv_1
xIinv[7] otrip_decoded_avdd[7] VGND VNB VPB VPWR otrip_decoded_b_avdd[7] sky130_fd_sc_hvl__inv_1
xIinv[6] otrip_decoded_avdd[6] VGND VNB VPB VPWR otrip_decoded_b_avdd[6] sky130_fd_sc_hvl__inv_1
xIinv[5] otrip_decoded_avdd[5] VGND VNB VPB VPWR otrip_decoded_b_avdd[5] sky130_fd_sc_hvl__inv_1
xIinv[4] otrip_decoded_avdd[4] VGND VNB VPB VPWR otrip_decoded_b_avdd[4] sky130_fd_sc_hvl__inv_1
xIinv[3] otrip_decoded_avdd[3] VGND VNB VPB VPWR otrip_decoded_b_avdd[3] sky130_fd_sc_hvl__inv_1
xIinv[2] otrip_decoded_avdd[2] VGND VNB VPB VPWR otrip_decoded_b_avdd[2] sky130_fd_sc_hvl__inv_1
xIinv[1] otrip_decoded_avdd[1] VGND VNB VPB VPWR otrip_decoded_b_avdd[1] sky130_fd_sc_hvl__inv_1
xIinv[0] otrip_decoded_avdd[0] VGND VNB VPB VPWR otrip_decoded_b_avdd[0] sky130_fd_sc_hvl__inv_1
.ends


* expanding   symbol:  comparator.sym # of pins=7
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/comparator.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/comparator.sch
.subckt comparator avdd ibias out ena vinn vinp avss
*.PININFO ena:I avdd:I avss:I ibias:I vinn:I vinp:I out:O
XMb vn vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMta vt vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMl0 vn ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMinv0 ena_b ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMinv1 ena_b ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMi0 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=4
XMi1 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=4
XMld1 vpp vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMh1 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1.5 nf=1 m=2
XMh0 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1.5 nf=1 m=2
XMld0 vnn vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMpp1 n0 vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMnn1 n0 vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMpp0 vm vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMnn0 vm vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMinv3 n1 n0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 nf=1 m=2
XMinv2 n1 n0 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 nf=1 m=2
XMinv5 out n1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 nf=1 m=8
XMinv4 out n1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 nf=1 m=8
XMl1 vm ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMl3 vnn ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMl4 vpp ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMt1 ibias ena vn avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMt0 vn ena_b ibias avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMl2 n0 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  ibias_gen.sym # of pins=8
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/ibias_gen.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__overvoltage/xschem/ibias_gen.sch
.subckt ibias_gen avdd itest ibias ibg_200n vbg_1v2 isrc_sel ena avss
*.PININFO vbg_1v2:I ena:I ibias:O ibg_200n:I isrc_sel:I avdd:I avss:I itest:O
XR1 avss net3 avss sky130_fd_pr__res_xhigh_po W=2 L=1000 mult=1 m=1
XQ1 avss avss net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XM17 net1 vbg_1v2 vn0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=10
XMt9 net1 ena_b net4 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMn0 vn0 vn0 net2 avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMp0 vn0 vp0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMn1 vp0 vn0 net3 avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMp1 vp0 vp0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMp ibias vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMt0 vp0 isrc_sel vp avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt1 vp isrc_sel_b vp0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMl6 vp ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl3 vp0 ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl1 vn0 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMnn1 vp1 vn1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 m=8
XMnn0 vn1 vn1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 m=2
XMl9 vn1 isrc_sel_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMt6 net5 isrc_sel vn1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt7 vn1 isrc_sel_b net6 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMpp1 vp1 vp1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMt2 vp isrc_sel_b vp1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt3 vp1 isrc_sel vp avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt4 ibg_200n ena net5 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt5 net6 ena_b ibg_200n avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMl7 vp1 isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl8 vp1 ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl10 vn1 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl2 vp0 isrc_sel_b avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl0 vn0 isrc_sel avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMt8 net4 isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMn2 ena_b ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMp2 ena_b ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMn3 isrc_sel_b isrc_sel avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMp3 isrc_sel_b isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMtst itest vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
.ends

.end
