magic
tech sky130A
magscale 1 2
timestamp 1712109191
<< error_p >>
rect -29 -129 29 129
<< pwell >>
rect -3515 -3194 3515 3194
<< mvnmos >>
rect -3287 1936 -1687 2936
rect -1629 1936 -29 2936
rect 29 1936 1629 2936
rect 1687 1936 3287 2936
rect -3287 718 -1687 1718
rect -1629 718 -29 1718
rect 29 718 1629 1718
rect 1687 718 3287 1718
rect -3287 -500 -1687 500
rect -1629 -500 -29 500
rect 29 -500 1629 500
rect 1687 -500 3287 500
rect -3287 -1718 -1687 -718
rect -1629 -1718 -29 -718
rect 29 -1718 1629 -718
rect 1687 -1718 3287 -718
rect -3287 -2936 -1687 -1936
rect -1629 -2936 -29 -1936
rect 29 -2936 1629 -1936
rect 1687 -2936 3287 -1936
<< mvndiff >>
rect -3345 2924 -3287 2936
rect -3345 1948 -3333 2924
rect -3299 1948 -3287 2924
rect -3345 1936 -3287 1948
rect -1687 2924 -1629 2936
rect -1687 1948 -1675 2924
rect -1641 1948 -1629 2924
rect -1687 1936 -1629 1948
rect -29 2924 29 2936
rect -29 1948 -17 2924
rect 17 1948 29 2924
rect -29 1936 29 1948
rect 1629 2924 1687 2936
rect 1629 1948 1641 2924
rect 1675 1948 1687 2924
rect 1629 1936 1687 1948
rect 3287 2924 3345 2936
rect 3287 1948 3299 2924
rect 3333 1948 3345 2924
rect 3287 1936 3345 1948
rect -3345 1706 -3287 1718
rect -3345 730 -3333 1706
rect -3299 730 -3287 1706
rect -3345 718 -3287 730
rect -1687 1706 -1629 1718
rect -1687 730 -1675 1706
rect -1641 730 -1629 1706
rect -1687 718 -1629 730
rect -29 1706 29 1718
rect -29 730 -17 1706
rect 17 730 29 1706
rect -29 718 29 730
rect 1629 1706 1687 1718
rect 1629 730 1641 1706
rect 1675 730 1687 1706
rect 1629 718 1687 730
rect 3287 1706 3345 1718
rect 3287 730 3299 1706
rect 3333 730 3345 1706
rect 3287 718 3345 730
rect -3345 488 -3287 500
rect -3345 -488 -3333 488
rect -3299 -488 -3287 488
rect -3345 -500 -3287 -488
rect -1687 488 -1629 500
rect -1687 -488 -1675 488
rect -1641 -488 -1629 488
rect -1687 -500 -1629 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 1629 488 1687 500
rect 1629 -488 1641 488
rect 1675 -488 1687 488
rect 1629 -500 1687 -488
rect 3287 488 3345 500
rect 3287 -488 3299 488
rect 3333 -488 3345 488
rect 3287 -500 3345 -488
rect -3345 -730 -3287 -718
rect -3345 -1706 -3333 -730
rect -3299 -1706 -3287 -730
rect -3345 -1718 -3287 -1706
rect -1687 -730 -1629 -718
rect -1687 -1706 -1675 -730
rect -1641 -1706 -1629 -730
rect -1687 -1718 -1629 -1706
rect -29 -730 29 -718
rect -29 -1706 -17 -730
rect 17 -1706 29 -730
rect -29 -1718 29 -1706
rect 1629 -730 1687 -718
rect 1629 -1706 1641 -730
rect 1675 -1706 1687 -730
rect 1629 -1718 1687 -1706
rect 3287 -730 3345 -718
rect 3287 -1706 3299 -730
rect 3333 -1706 3345 -730
rect 3287 -1718 3345 -1706
rect -3345 -1948 -3287 -1936
rect -3345 -2924 -3333 -1948
rect -3299 -2924 -3287 -1948
rect -3345 -2936 -3287 -2924
rect -1687 -1948 -1629 -1936
rect -1687 -2924 -1675 -1948
rect -1641 -2924 -1629 -1948
rect -1687 -2936 -1629 -2924
rect -29 -1948 29 -1936
rect -29 -2924 -17 -1948
rect 17 -2924 29 -1948
rect -29 -2936 29 -2924
rect 1629 -1948 1687 -1936
rect 1629 -2924 1641 -1948
rect 1675 -2924 1687 -1948
rect 1629 -2936 1687 -2924
rect 3287 -1948 3345 -1936
rect 3287 -2924 3299 -1948
rect 3333 -2924 3345 -1948
rect 3287 -2936 3345 -2924
<< mvndiffc >>
rect -3333 1948 -3299 2924
rect -1675 1948 -1641 2924
rect -17 1948 17 2924
rect 1641 1948 1675 2924
rect 3299 1948 3333 2924
rect -3333 730 -3299 1706
rect -1675 730 -1641 1706
rect -17 730 17 1706
rect 1641 730 1675 1706
rect 3299 730 3333 1706
rect -3333 -488 -3299 488
rect -1675 -488 -1641 488
rect -17 -488 17 488
rect 1641 -488 1675 488
rect 3299 -488 3333 488
rect -3333 -1706 -3299 -730
rect -1675 -1706 -1641 -730
rect -17 -1706 17 -730
rect 1641 -1706 1675 -730
rect 3299 -1706 3333 -730
rect -3333 -2924 -3299 -1948
rect -1675 -2924 -1641 -1948
rect -17 -2924 17 -1948
rect 1641 -2924 1675 -1948
rect 3299 -2924 3333 -1948
<< mvpsubdiff >>
rect -3479 3146 3479 3158
rect -3479 3112 -3371 3146
rect 3371 3112 3479 3146
rect -3479 3100 3479 3112
rect -3479 3050 -3421 3100
rect -3479 -3050 -3467 3050
rect -3433 -3050 -3421 3050
rect 3421 3050 3479 3100
rect -3479 -3100 -3421 -3050
rect 3421 -3050 3433 3050
rect 3467 -3050 3479 3050
rect 3421 -3100 3479 -3050
rect -3479 -3112 3479 -3100
rect -3479 -3146 -3371 -3112
rect 3371 -3146 3479 -3112
rect -3479 -3158 3479 -3146
<< mvpsubdiffcont >>
rect -3371 3112 3371 3146
rect -3467 -3050 -3433 3050
rect 3433 -3050 3467 3050
rect -3371 -3146 3371 -3112
<< poly >>
rect -3287 3008 -1687 3024
rect -3287 2974 -3271 3008
rect -1703 2974 -1687 3008
rect -3287 2936 -1687 2974
rect -1629 3008 -29 3024
rect -1629 2974 -1613 3008
rect -45 2974 -29 3008
rect -1629 2936 -29 2974
rect 29 3008 1629 3024
rect 29 2974 45 3008
rect 1613 2974 1629 3008
rect 29 2936 1629 2974
rect 1687 3008 3287 3024
rect 1687 2974 1703 3008
rect 3271 2974 3287 3008
rect 1687 2936 3287 2974
rect -3287 1898 -1687 1936
rect -3287 1864 -3271 1898
rect -1703 1864 -1687 1898
rect -3287 1848 -1687 1864
rect -1629 1898 -29 1936
rect -1629 1864 -1613 1898
rect -45 1864 -29 1898
rect -1629 1848 -29 1864
rect 29 1898 1629 1936
rect 29 1864 45 1898
rect 1613 1864 1629 1898
rect 29 1848 1629 1864
rect 1687 1898 3287 1936
rect 1687 1864 1703 1898
rect 3271 1864 3287 1898
rect 1687 1848 3287 1864
rect -3287 1790 -1687 1806
rect -3287 1756 -3271 1790
rect -1703 1756 -1687 1790
rect -3287 1718 -1687 1756
rect -1629 1790 -29 1806
rect -1629 1756 -1613 1790
rect -45 1756 -29 1790
rect -1629 1718 -29 1756
rect 29 1790 1629 1806
rect 29 1756 45 1790
rect 1613 1756 1629 1790
rect 29 1718 1629 1756
rect 1687 1790 3287 1806
rect 1687 1756 1703 1790
rect 3271 1756 3287 1790
rect 1687 1718 3287 1756
rect -3287 680 -1687 718
rect -3287 646 -3271 680
rect -1703 646 -1687 680
rect -3287 630 -1687 646
rect -1629 680 -29 718
rect -1629 646 -1613 680
rect -45 646 -29 680
rect -1629 630 -29 646
rect 29 680 1629 718
rect 29 646 45 680
rect 1613 646 1629 680
rect 29 630 1629 646
rect 1687 680 3287 718
rect 1687 646 1703 680
rect 3271 646 3287 680
rect 1687 630 3287 646
rect -3287 572 -1687 588
rect -3287 538 -3271 572
rect -1703 538 -1687 572
rect -3287 500 -1687 538
rect -1629 572 -29 588
rect -1629 538 -1613 572
rect -45 538 -29 572
rect -1629 500 -29 538
rect 29 572 1629 588
rect 29 538 45 572
rect 1613 538 1629 572
rect 29 500 1629 538
rect 1687 572 3287 588
rect 1687 538 1703 572
rect 3271 538 3287 572
rect 1687 500 3287 538
rect -3287 -538 -1687 -500
rect -3287 -572 -3271 -538
rect -1703 -572 -1687 -538
rect -3287 -588 -1687 -572
rect -1629 -538 -29 -500
rect -1629 -572 -1613 -538
rect -45 -572 -29 -538
rect -1629 -588 -29 -572
rect 29 -538 1629 -500
rect 29 -572 45 -538
rect 1613 -572 1629 -538
rect 29 -588 1629 -572
rect 1687 -538 3287 -500
rect 1687 -572 1703 -538
rect 3271 -572 3287 -538
rect 1687 -588 3287 -572
rect -3287 -646 -1687 -630
rect -3287 -680 -3271 -646
rect -1703 -680 -1687 -646
rect -3287 -718 -1687 -680
rect -1629 -646 -29 -630
rect -1629 -680 -1613 -646
rect -45 -680 -29 -646
rect -1629 -718 -29 -680
rect 29 -646 1629 -630
rect 29 -680 45 -646
rect 1613 -680 1629 -646
rect 29 -718 1629 -680
rect 1687 -646 3287 -630
rect 1687 -680 1703 -646
rect 3271 -680 3287 -646
rect 1687 -718 3287 -680
rect -3287 -1756 -1687 -1718
rect -3287 -1790 -3271 -1756
rect -1703 -1790 -1687 -1756
rect -3287 -1806 -1687 -1790
rect -1629 -1756 -29 -1718
rect -1629 -1790 -1613 -1756
rect -45 -1790 -29 -1756
rect -1629 -1806 -29 -1790
rect 29 -1756 1629 -1718
rect 29 -1790 45 -1756
rect 1613 -1790 1629 -1756
rect 29 -1806 1629 -1790
rect 1687 -1756 3287 -1718
rect 1687 -1790 1703 -1756
rect 3271 -1790 3287 -1756
rect 1687 -1806 3287 -1790
rect -3287 -1864 -1687 -1848
rect -3287 -1898 -3271 -1864
rect -1703 -1898 -1687 -1864
rect -3287 -1936 -1687 -1898
rect -1629 -1864 -29 -1848
rect -1629 -1898 -1613 -1864
rect -45 -1898 -29 -1864
rect -1629 -1936 -29 -1898
rect 29 -1864 1629 -1848
rect 29 -1898 45 -1864
rect 1613 -1898 1629 -1864
rect 29 -1936 1629 -1898
rect 1687 -1864 3287 -1848
rect 1687 -1898 1703 -1864
rect 3271 -1898 3287 -1864
rect 1687 -1936 3287 -1898
rect -3287 -2974 -1687 -2936
rect -3287 -3008 -3271 -2974
rect -1703 -3008 -1687 -2974
rect -3287 -3024 -1687 -3008
rect -1629 -2974 -29 -2936
rect -1629 -3008 -1613 -2974
rect -45 -3008 -29 -2974
rect -1629 -3024 -29 -3008
rect 29 -2974 1629 -2936
rect 29 -3008 45 -2974
rect 1613 -3008 1629 -2974
rect 29 -3024 1629 -3008
rect 1687 -2974 3287 -2936
rect 1687 -3008 1703 -2974
rect 3271 -3008 3287 -2974
rect 1687 -3024 3287 -3008
<< polycont >>
rect -3271 2974 -1703 3008
rect -1613 2974 -45 3008
rect 45 2974 1613 3008
rect 1703 2974 3271 3008
rect -3271 1864 -1703 1898
rect -1613 1864 -45 1898
rect 45 1864 1613 1898
rect 1703 1864 3271 1898
rect -3271 1756 -1703 1790
rect -1613 1756 -45 1790
rect 45 1756 1613 1790
rect 1703 1756 3271 1790
rect -3271 646 -1703 680
rect -1613 646 -45 680
rect 45 646 1613 680
rect 1703 646 3271 680
rect -3271 538 -1703 572
rect -1613 538 -45 572
rect 45 538 1613 572
rect 1703 538 3271 572
rect -3271 -572 -1703 -538
rect -1613 -572 -45 -538
rect 45 -572 1613 -538
rect 1703 -572 3271 -538
rect -3271 -680 -1703 -646
rect -1613 -680 -45 -646
rect 45 -680 1613 -646
rect 1703 -680 3271 -646
rect -3271 -1790 -1703 -1756
rect -1613 -1790 -45 -1756
rect 45 -1790 1613 -1756
rect 1703 -1790 3271 -1756
rect -3271 -1898 -1703 -1864
rect -1613 -1898 -45 -1864
rect 45 -1898 1613 -1864
rect 1703 -1898 3271 -1864
rect -3271 -3008 -1703 -2974
rect -1613 -3008 -45 -2974
rect 45 -3008 1613 -2974
rect 1703 -3008 3271 -2974
<< locali >>
rect -3467 3112 -3371 3146
rect 3371 3112 3467 3146
rect -3467 3050 -3433 3112
rect 3433 3050 3467 3112
rect -3287 2974 -3271 3008
rect -1703 2974 -1687 3008
rect -1629 2974 -1613 3008
rect -45 2974 -29 3008
rect 29 2974 45 3008
rect 1613 2974 1629 3008
rect 1687 2974 1703 3008
rect 3271 2974 3287 3008
rect -3333 2924 -3299 2940
rect -3333 1932 -3299 1948
rect -1675 2924 -1641 2940
rect -1675 1932 -1641 1948
rect -17 2924 17 2940
rect -17 1932 17 1948
rect 1641 2924 1675 2940
rect 1641 1932 1675 1948
rect 3299 2924 3333 2940
rect 3299 1932 3333 1948
rect -3287 1864 -3271 1898
rect -1703 1864 -1687 1898
rect -1629 1864 -1613 1898
rect -45 1864 -29 1898
rect 29 1864 45 1898
rect 1613 1864 1629 1898
rect 1687 1864 1703 1898
rect 3271 1864 3287 1898
rect -3287 1756 -3271 1790
rect -1703 1756 -1687 1790
rect -1629 1756 -1613 1790
rect -45 1756 -29 1790
rect 29 1756 45 1790
rect 1613 1756 1629 1790
rect 1687 1756 1703 1790
rect 3271 1756 3287 1790
rect -3333 1706 -3299 1722
rect -3333 714 -3299 730
rect -1675 1706 -1641 1722
rect -1675 714 -1641 730
rect -17 1706 17 1722
rect -17 714 17 730
rect 1641 1706 1675 1722
rect 1641 714 1675 730
rect 3299 1706 3333 1722
rect 3299 714 3333 730
rect -3287 646 -3271 680
rect -1703 646 -1687 680
rect -1629 646 -1613 680
rect -45 646 -29 680
rect 29 646 45 680
rect 1613 646 1629 680
rect 1687 646 1703 680
rect 3271 646 3287 680
rect -3287 538 -3271 572
rect -1703 538 -1687 572
rect -1629 538 -1613 572
rect -45 538 -29 572
rect 29 538 45 572
rect 1613 538 1629 572
rect 1687 538 1703 572
rect 3271 538 3287 572
rect -3333 488 -3299 504
rect -3333 -504 -3299 -488
rect -1675 488 -1641 504
rect -1675 -504 -1641 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 1641 488 1675 504
rect 1641 -504 1675 -488
rect 3299 488 3333 504
rect 3299 -504 3333 -488
rect -3287 -572 -3271 -538
rect -1703 -572 -1687 -538
rect -1629 -572 -1613 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 1613 -572 1629 -538
rect 1687 -572 1703 -538
rect 3271 -572 3287 -538
rect -3287 -680 -3271 -646
rect -1703 -680 -1687 -646
rect -1629 -680 -1613 -646
rect -45 -680 -29 -646
rect 29 -680 45 -646
rect 1613 -680 1629 -646
rect 1687 -680 1703 -646
rect 3271 -680 3287 -646
rect -3333 -730 -3299 -714
rect -3333 -1722 -3299 -1706
rect -1675 -730 -1641 -714
rect -1675 -1722 -1641 -1706
rect -17 -730 17 -714
rect -17 -1722 17 -1706
rect 1641 -730 1675 -714
rect 1641 -1722 1675 -1706
rect 3299 -730 3333 -714
rect 3299 -1722 3333 -1706
rect -3287 -1790 -3271 -1756
rect -1703 -1790 -1687 -1756
rect -1629 -1790 -1613 -1756
rect -45 -1790 -29 -1756
rect 29 -1790 45 -1756
rect 1613 -1790 1629 -1756
rect 1687 -1790 1703 -1756
rect 3271 -1790 3287 -1756
rect -3287 -1898 -3271 -1864
rect -1703 -1898 -1687 -1864
rect -1629 -1898 -1613 -1864
rect -45 -1898 -29 -1864
rect 29 -1898 45 -1864
rect 1613 -1898 1629 -1864
rect 1687 -1898 1703 -1864
rect 3271 -1898 3287 -1864
rect -3333 -1948 -3299 -1932
rect -3333 -2940 -3299 -2924
rect -1675 -1948 -1641 -1932
rect -1675 -2940 -1641 -2924
rect -17 -1948 17 -1932
rect -17 -2940 17 -2924
rect 1641 -1948 1675 -1932
rect 1641 -2940 1675 -2924
rect 3299 -1948 3333 -1932
rect 3299 -2940 3333 -2924
rect -3287 -3008 -3271 -2974
rect -1703 -3008 -1687 -2974
rect -1629 -3008 -1613 -2974
rect -45 -3008 -29 -2974
rect 29 -3008 45 -2974
rect 1613 -3008 1629 -2974
rect 1687 -3008 1703 -2974
rect 3271 -3008 3287 -2974
rect -3467 -3112 -3433 -3050
rect 3433 -3112 3467 -3050
rect -3467 -3146 -3371 -3112
rect 3371 -3146 3467 -3112
<< viali >>
rect -3271 2974 -1703 3008
rect -1613 2974 -45 3008
rect 45 2974 1613 3008
rect 1703 2974 3271 3008
rect -3333 1948 -3299 2924
rect -1675 1948 -1641 2924
rect -17 1948 17 2924
rect 1641 1948 1675 2924
rect 3299 1948 3333 2924
rect -3271 1864 -1703 1898
rect -1613 1864 -45 1898
rect 45 1864 1613 1898
rect 1703 1864 3271 1898
rect -3271 1756 -1703 1790
rect -1613 1756 -45 1790
rect 45 1756 1613 1790
rect 1703 1756 3271 1790
rect -3333 730 -3299 1706
rect -1675 730 -1641 1706
rect -17 730 17 1706
rect 1641 730 1675 1706
rect 3299 730 3333 1706
rect -3271 646 -1703 680
rect -1613 646 -45 680
rect 45 646 1613 680
rect 1703 646 3271 680
rect -3271 538 -1703 572
rect -1613 538 -45 572
rect 45 538 1613 572
rect 1703 538 3271 572
rect -3333 -488 -3299 488
rect -1675 -488 -1641 488
rect -17 -488 17 488
rect 1641 -488 1675 488
rect 3299 -488 3333 488
rect -3271 -572 -1703 -538
rect -1613 -572 -45 -538
rect 45 -572 1613 -538
rect 1703 -572 3271 -538
rect -3271 -680 -1703 -646
rect -1613 -680 -45 -646
rect 45 -680 1613 -646
rect 1703 -680 3271 -646
rect -3333 -1706 -3299 -730
rect -1675 -1706 -1641 -730
rect -17 -1706 17 -730
rect 1641 -1706 1675 -730
rect 3299 -1706 3333 -730
rect -3271 -1790 -1703 -1756
rect -1613 -1790 -45 -1756
rect 45 -1790 1613 -1756
rect 1703 -1790 3271 -1756
rect -3271 -1898 -1703 -1864
rect -1613 -1898 -45 -1864
rect 45 -1898 1613 -1864
rect 1703 -1898 3271 -1864
rect -3333 -2924 -3299 -1948
rect -1675 -2924 -1641 -1948
rect -17 -2924 17 -1948
rect 1641 -2924 1675 -1948
rect 3299 -2924 3333 -1948
rect -3271 -3008 -1703 -2974
rect -1613 -3008 -45 -2974
rect 45 -3008 1613 -2974
rect 1703 -3008 3271 -2974
<< metal1 >>
rect -3283 3008 -1691 3014
rect -3283 2974 -3271 3008
rect -1703 2974 -1691 3008
rect -3283 2968 -1691 2974
rect -1625 3008 -33 3014
rect -1625 2974 -1613 3008
rect -45 2974 -33 3008
rect -1625 2968 -33 2974
rect 33 3008 1625 3014
rect 33 2974 45 3008
rect 1613 2974 1625 3008
rect 33 2968 1625 2974
rect 1691 3008 3283 3014
rect 1691 2974 1703 3008
rect 3271 2974 3283 3008
rect 1691 2968 3283 2974
rect -3339 2924 -3293 2936
rect -3339 1948 -3333 2924
rect -3299 1948 -3293 2924
rect -3339 1936 -3293 1948
rect -1681 2924 -1635 2936
rect -1681 1948 -1675 2924
rect -1641 1948 -1635 2924
rect -1681 1936 -1635 1948
rect -23 2924 23 2936
rect -23 1948 -17 2924
rect 17 1948 23 2924
rect -23 1936 23 1948
rect 1635 2924 1681 2936
rect 1635 1948 1641 2924
rect 1675 1948 1681 2924
rect 1635 1936 1681 1948
rect 3293 2924 3339 2936
rect 3293 1948 3299 2924
rect 3333 1948 3339 2924
rect 3293 1936 3339 1948
rect -3283 1898 -1691 1904
rect -3283 1864 -3271 1898
rect -1703 1864 -1691 1898
rect -3283 1858 -1691 1864
rect -1625 1898 -33 1904
rect -1625 1864 -1613 1898
rect -45 1864 -33 1898
rect -1625 1858 -33 1864
rect 33 1898 1625 1904
rect 33 1864 45 1898
rect 1613 1864 1625 1898
rect 33 1858 1625 1864
rect 1691 1898 3283 1904
rect 1691 1864 1703 1898
rect 3271 1864 3283 1898
rect 1691 1858 3283 1864
rect -3283 1790 -1691 1796
rect -3283 1756 -3271 1790
rect -1703 1756 -1691 1790
rect -3283 1750 -1691 1756
rect -1625 1790 -33 1796
rect -1625 1756 -1613 1790
rect -45 1756 -33 1790
rect -1625 1750 -33 1756
rect 33 1790 1625 1796
rect 33 1756 45 1790
rect 1613 1756 1625 1790
rect 33 1750 1625 1756
rect 1691 1790 3283 1796
rect 1691 1756 1703 1790
rect 3271 1756 3283 1790
rect 1691 1750 3283 1756
rect -3339 1706 -3293 1718
rect -3339 730 -3333 1706
rect -3299 730 -3293 1706
rect -3339 718 -3293 730
rect -1681 1706 -1635 1718
rect -1681 730 -1675 1706
rect -1641 730 -1635 1706
rect -1681 718 -1635 730
rect -23 1706 23 1718
rect -23 730 -17 1706
rect 17 730 23 1706
rect -23 718 23 730
rect 1635 1706 1681 1718
rect 1635 730 1641 1706
rect 1675 730 1681 1706
rect 1635 718 1681 730
rect 3293 1706 3339 1718
rect 3293 730 3299 1706
rect 3333 730 3339 1706
rect 3293 718 3339 730
rect -3283 680 -1691 686
rect -3283 646 -3271 680
rect -1703 646 -1691 680
rect -3283 640 -1691 646
rect -1625 680 -33 686
rect -1625 646 -1613 680
rect -45 646 -33 680
rect -1625 640 -33 646
rect 33 680 1625 686
rect 33 646 45 680
rect 1613 646 1625 680
rect 33 640 1625 646
rect 1691 680 3283 686
rect 1691 646 1703 680
rect 3271 646 3283 680
rect 1691 640 3283 646
rect -3283 572 -1691 578
rect -3283 538 -3271 572
rect -1703 538 -1691 572
rect -3283 532 -1691 538
rect -1625 572 -33 578
rect -1625 538 -1613 572
rect -45 538 -33 572
rect -1625 532 -33 538
rect 33 572 1625 578
rect 33 538 45 572
rect 1613 538 1625 572
rect 33 532 1625 538
rect 1691 572 3283 578
rect 1691 538 1703 572
rect 3271 538 3283 572
rect 1691 532 3283 538
rect -3339 488 -3293 500
rect -3339 -488 -3333 488
rect -3299 -488 -3293 488
rect -3339 -500 -3293 -488
rect -1681 488 -1635 500
rect -1681 -488 -1675 488
rect -1641 -488 -1635 488
rect -1681 -500 -1635 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 1635 488 1681 500
rect 1635 -488 1641 488
rect 1675 -488 1681 488
rect 1635 -500 1681 -488
rect 3293 488 3339 500
rect 3293 -488 3299 488
rect 3333 -488 3339 488
rect 3293 -500 3339 -488
rect -3283 -538 -1691 -532
rect -3283 -572 -3271 -538
rect -1703 -572 -1691 -538
rect -3283 -578 -1691 -572
rect -1625 -538 -33 -532
rect -1625 -572 -1613 -538
rect -45 -572 -33 -538
rect -1625 -578 -33 -572
rect 33 -538 1625 -532
rect 33 -572 45 -538
rect 1613 -572 1625 -538
rect 33 -578 1625 -572
rect 1691 -538 3283 -532
rect 1691 -572 1703 -538
rect 3271 -572 3283 -538
rect 1691 -578 3283 -572
rect -3283 -646 -1691 -640
rect -3283 -680 -3271 -646
rect -1703 -680 -1691 -646
rect -3283 -686 -1691 -680
rect -1625 -646 -33 -640
rect -1625 -680 -1613 -646
rect -45 -680 -33 -646
rect -1625 -686 -33 -680
rect 33 -646 1625 -640
rect 33 -680 45 -646
rect 1613 -680 1625 -646
rect 33 -686 1625 -680
rect 1691 -646 3283 -640
rect 1691 -680 1703 -646
rect 3271 -680 3283 -646
rect 1691 -686 3283 -680
rect -3339 -730 -3293 -718
rect -3339 -1706 -3333 -730
rect -3299 -1706 -3293 -730
rect -3339 -1718 -3293 -1706
rect -1681 -730 -1635 -718
rect -1681 -1706 -1675 -730
rect -1641 -1706 -1635 -730
rect -1681 -1718 -1635 -1706
rect -23 -730 23 -718
rect -23 -1706 -17 -730
rect 17 -1706 23 -730
rect -23 -1718 23 -1706
rect 1635 -730 1681 -718
rect 1635 -1706 1641 -730
rect 1675 -1706 1681 -730
rect 1635 -1718 1681 -1706
rect 3293 -730 3339 -718
rect 3293 -1706 3299 -730
rect 3333 -1706 3339 -730
rect 3293 -1718 3339 -1706
rect -3283 -1756 -1691 -1750
rect -3283 -1790 -3271 -1756
rect -1703 -1790 -1691 -1756
rect -3283 -1796 -1691 -1790
rect -1625 -1756 -33 -1750
rect -1625 -1790 -1613 -1756
rect -45 -1790 -33 -1756
rect -1625 -1796 -33 -1790
rect 33 -1756 1625 -1750
rect 33 -1790 45 -1756
rect 1613 -1790 1625 -1756
rect 33 -1796 1625 -1790
rect 1691 -1756 3283 -1750
rect 1691 -1790 1703 -1756
rect 3271 -1790 3283 -1756
rect 1691 -1796 3283 -1790
rect -3283 -1864 -1691 -1858
rect -3283 -1898 -3271 -1864
rect -1703 -1898 -1691 -1864
rect -3283 -1904 -1691 -1898
rect -1625 -1864 -33 -1858
rect -1625 -1898 -1613 -1864
rect -45 -1898 -33 -1864
rect -1625 -1904 -33 -1898
rect 33 -1864 1625 -1858
rect 33 -1898 45 -1864
rect 1613 -1898 1625 -1864
rect 33 -1904 1625 -1898
rect 1691 -1864 3283 -1858
rect 1691 -1898 1703 -1864
rect 3271 -1898 3283 -1864
rect 1691 -1904 3283 -1898
rect -3339 -1948 -3293 -1936
rect -3339 -2924 -3333 -1948
rect -3299 -2924 -3293 -1948
rect -3339 -2936 -3293 -2924
rect -1681 -1948 -1635 -1936
rect -1681 -2924 -1675 -1948
rect -1641 -2924 -1635 -1948
rect -1681 -2936 -1635 -2924
rect -23 -1948 23 -1936
rect -23 -2924 -17 -1948
rect 17 -2924 23 -1948
rect -23 -2936 23 -2924
rect 1635 -1948 1681 -1936
rect 1635 -2924 1641 -1948
rect 1675 -2924 1681 -1948
rect 1635 -2936 1681 -2924
rect 3293 -1948 3339 -1936
rect 3293 -2924 3299 -1948
rect 3333 -2924 3339 -1948
rect 3293 -2936 3339 -2924
rect -3283 -2974 -1691 -2968
rect -3283 -3008 -3271 -2974
rect -1703 -3008 -1691 -2974
rect -3283 -3014 -1691 -3008
rect -1625 -2974 -33 -2968
rect -1625 -3008 -1613 -2974
rect -45 -3008 -33 -2974
rect -1625 -3014 -33 -3008
rect 33 -2974 1625 -2968
rect 33 -3008 45 -2974
rect 1613 -3008 1625 -2974
rect 33 -3014 1625 -3008
rect 1691 -2974 3283 -2968
rect 1691 -3008 1703 -2974
rect 3271 -3008 3283 -2974
rect 1691 -3014 3283 -3008
<< properties >>
string FIXED_BBOX -3450 -3129 3450 3129
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 8 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
