magic
tech sky130A
magscale 1 2
timestamp 1712457293
<< metal3 >>
rect -3186 9332 3186 9360
rect -3186 3308 3102 9332
rect 3166 3308 3186 9332
rect -3186 3280 3186 3308
rect -3186 3012 3186 3040
rect -3186 -3012 3102 3012
rect 3166 -3012 3186 3012
rect -3186 -3040 3186 -3012
rect -3186 -3308 3186 -3280
rect -3186 -9332 3102 -3308
rect 3166 -9332 3186 -3308
rect -3186 -9360 3186 -9332
<< via3 >>
rect 3102 3308 3166 9332
rect 3102 -3012 3166 3012
rect 3102 -9332 3166 -3308
<< mimcap >>
rect -3146 9280 2854 9320
rect -3146 3360 -3106 9280
rect 2814 3360 2854 9280
rect -3146 3320 2854 3360
rect -3146 2960 2854 3000
rect -3146 -2960 -3106 2960
rect 2814 -2960 2854 2960
rect -3146 -3000 2854 -2960
rect -3146 -3360 2854 -3320
rect -3146 -9280 -3106 -3360
rect 2814 -9280 2854 -3360
rect -3146 -9320 2854 -9280
<< mimcapcontact >>
rect -3106 3360 2814 9280
rect -3106 -2960 2814 2960
rect -3106 -9280 2814 -3360
<< metal4 >>
rect -198 9281 -94 9480
rect 3082 9332 3186 9480
rect -3107 9280 2815 9281
rect -3107 3360 -3106 9280
rect 2814 3360 2815 9280
rect -3107 3359 2815 3360
rect -198 2961 -94 3359
rect 3082 3308 3102 9332
rect 3166 3308 3186 9332
rect 3082 3012 3186 3308
rect -3107 2960 2815 2961
rect -3107 -2960 -3106 2960
rect 2814 -2960 2815 2960
rect -3107 -2961 2815 -2960
rect -198 -3359 -94 -2961
rect 3082 -3012 3102 3012
rect 3166 -3012 3186 3012
rect 3082 -3308 3186 -3012
rect -3107 -3360 2815 -3359
rect -3107 -9280 -3106 -3360
rect 2814 -9280 2815 -3360
rect -3107 -9281 2815 -9280
rect -198 -9480 -94 -9281
rect 3082 -9332 3102 -3308
rect 3166 -9332 3186 -3308
rect 3082 -9480 3186 -9332
<< properties >>
string FIXED_BBOX -3186 3280 2894 9360
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
