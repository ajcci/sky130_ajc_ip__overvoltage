magic
tech sky130A
timestamp 1711636687
<< nwell >>
rect -4259 -249 4259 249
<< mvpmos >>
rect -4130 59 -3330 101
rect -3301 59 -2501 101
rect -2472 59 -1672 101
rect -1643 59 -843 101
rect -814 59 -14 101
rect 14 59 814 101
rect 843 59 1643 101
rect 1672 59 2472 101
rect 2501 59 3301 101
rect 3330 59 4130 101
rect -4130 -101 -3330 -59
rect -3301 -101 -2501 -59
rect -2472 -101 -1672 -59
rect -1643 -101 -843 -59
rect -814 -101 -14 -59
rect 14 -101 814 -59
rect 843 -101 1643 -59
rect 1672 -101 2472 -59
rect 2501 -101 3301 -59
rect 3330 -101 4130 -59
<< mvpdiff >>
rect -4159 95 -4130 101
rect -4159 65 -4153 95
rect -4136 65 -4130 95
rect -4159 59 -4130 65
rect -3330 95 -3301 101
rect -3330 65 -3324 95
rect -3307 65 -3301 95
rect -3330 59 -3301 65
rect -2501 95 -2472 101
rect -2501 65 -2495 95
rect -2478 65 -2472 95
rect -2501 59 -2472 65
rect -1672 95 -1643 101
rect -1672 65 -1666 95
rect -1649 65 -1643 95
rect -1672 59 -1643 65
rect -843 95 -814 101
rect -843 65 -837 95
rect -820 65 -814 95
rect -843 59 -814 65
rect -14 95 14 101
rect -14 65 -8 95
rect 8 65 14 95
rect -14 59 14 65
rect 814 95 843 101
rect 814 65 820 95
rect 837 65 843 95
rect 814 59 843 65
rect 1643 95 1672 101
rect 1643 65 1649 95
rect 1666 65 1672 95
rect 1643 59 1672 65
rect 2472 95 2501 101
rect 2472 65 2478 95
rect 2495 65 2501 95
rect 2472 59 2501 65
rect 3301 95 3330 101
rect 3301 65 3307 95
rect 3324 65 3330 95
rect 3301 59 3330 65
rect 4130 95 4159 101
rect 4130 65 4136 95
rect 4153 65 4159 95
rect 4130 59 4159 65
rect -4159 -65 -4130 -59
rect -4159 -95 -4153 -65
rect -4136 -95 -4130 -65
rect -4159 -101 -4130 -95
rect -3330 -65 -3301 -59
rect -3330 -95 -3324 -65
rect -3307 -95 -3301 -65
rect -3330 -101 -3301 -95
rect -2501 -65 -2472 -59
rect -2501 -95 -2495 -65
rect -2478 -95 -2472 -65
rect -2501 -101 -2472 -95
rect -1672 -65 -1643 -59
rect -1672 -95 -1666 -65
rect -1649 -95 -1643 -65
rect -1672 -101 -1643 -95
rect -843 -65 -814 -59
rect -843 -95 -837 -65
rect -820 -95 -814 -65
rect -843 -101 -814 -95
rect -14 -65 14 -59
rect -14 -95 -8 -65
rect 8 -95 14 -65
rect -14 -101 14 -95
rect 814 -65 843 -59
rect 814 -95 820 -65
rect 837 -95 843 -65
rect 814 -101 843 -95
rect 1643 -65 1672 -59
rect 1643 -95 1649 -65
rect 1666 -95 1672 -65
rect 1643 -101 1672 -95
rect 2472 -65 2501 -59
rect 2472 -95 2478 -65
rect 2495 -95 2501 -65
rect 2472 -101 2501 -95
rect 3301 -65 3330 -59
rect 3301 -95 3307 -65
rect 3324 -95 3330 -65
rect 3301 -101 3330 -95
rect 4130 -65 4159 -59
rect 4130 -95 4136 -65
rect 4153 -95 4159 -65
rect 4130 -101 4159 -95
<< mvpdiffc >>
rect -4153 65 -4136 95
rect -3324 65 -3307 95
rect -2495 65 -2478 95
rect -1666 65 -1649 95
rect -837 65 -820 95
rect -8 65 8 95
rect 820 65 837 95
rect 1649 65 1666 95
rect 2478 65 2495 95
rect 3307 65 3324 95
rect 4136 65 4153 95
rect -4153 -95 -4136 -65
rect -3324 -95 -3307 -65
rect -2495 -95 -2478 -65
rect -1666 -95 -1649 -65
rect -837 -95 -820 -65
rect -8 -95 8 -65
rect 820 -95 837 -65
rect 1649 -95 1666 -65
rect 2478 -95 2495 -65
rect 3307 -95 3324 -65
rect 4136 -95 4153 -65
<< mvnsubdiff >>
rect -4226 210 4226 216
rect -4226 193 -4172 210
rect 4172 193 4226 210
rect -4226 187 4226 193
rect -4226 162 -4197 187
rect -4226 -162 -4220 162
rect -4203 -162 -4197 162
rect 4197 162 4226 187
rect -4226 -187 -4197 -162
rect 4197 -162 4203 162
rect 4220 -162 4226 162
rect 4197 -187 4226 -162
rect -4226 -193 4226 -187
rect -4226 -210 -4172 -193
rect 4172 -210 4226 -193
rect -4226 -216 4226 -210
<< mvnsubdiffcont >>
rect -4172 193 4172 210
rect -4220 -162 -4203 162
rect 4203 -162 4220 162
rect -4172 -210 4172 -193
<< poly >>
rect -4130 141 -3330 149
rect -4130 124 -4122 141
rect -3338 124 -3330 141
rect -4130 101 -3330 124
rect -3301 141 -2501 149
rect -3301 124 -3293 141
rect -2509 124 -2501 141
rect -3301 101 -2501 124
rect -2472 141 -1672 149
rect -2472 124 -2464 141
rect -1680 124 -1672 141
rect -2472 101 -1672 124
rect -1643 141 -843 149
rect -1643 124 -1635 141
rect -851 124 -843 141
rect -1643 101 -843 124
rect -814 141 -14 149
rect -814 124 -806 141
rect -22 124 -14 141
rect -814 101 -14 124
rect 14 141 814 149
rect 14 124 22 141
rect 806 124 814 141
rect 14 101 814 124
rect 843 141 1643 149
rect 843 124 851 141
rect 1635 124 1643 141
rect 843 101 1643 124
rect 1672 141 2472 149
rect 1672 124 1680 141
rect 2464 124 2472 141
rect 1672 101 2472 124
rect 2501 141 3301 149
rect 2501 124 2509 141
rect 3293 124 3301 141
rect 2501 101 3301 124
rect 3330 141 4130 149
rect 3330 124 3338 141
rect 4122 124 4130 141
rect 3330 101 4130 124
rect -4130 35 -3330 59
rect -4130 18 -4122 35
rect -3338 18 -3330 35
rect -4130 10 -3330 18
rect -3301 35 -2501 59
rect -3301 18 -3293 35
rect -2509 18 -2501 35
rect -3301 10 -2501 18
rect -2472 35 -1672 59
rect -2472 18 -2464 35
rect -1680 18 -1672 35
rect -2472 10 -1672 18
rect -1643 35 -843 59
rect -1643 18 -1635 35
rect -851 18 -843 35
rect -1643 10 -843 18
rect -814 35 -14 59
rect -814 18 -806 35
rect -22 18 -14 35
rect -814 10 -14 18
rect 14 35 814 59
rect 14 18 22 35
rect 806 18 814 35
rect 14 10 814 18
rect 843 35 1643 59
rect 843 18 851 35
rect 1635 18 1643 35
rect 843 10 1643 18
rect 1672 35 2472 59
rect 1672 18 1680 35
rect 2464 18 2472 35
rect 1672 10 2472 18
rect 2501 35 3301 59
rect 2501 18 2509 35
rect 3293 18 3301 35
rect 2501 10 3301 18
rect 3330 35 4130 59
rect 3330 18 3338 35
rect 4122 18 4130 35
rect 3330 10 4130 18
rect -4130 -18 -3330 -10
rect -4130 -35 -4122 -18
rect -3338 -35 -3330 -18
rect -4130 -59 -3330 -35
rect -3301 -18 -2501 -10
rect -3301 -35 -3293 -18
rect -2509 -35 -2501 -18
rect -3301 -59 -2501 -35
rect -2472 -18 -1672 -10
rect -2472 -35 -2464 -18
rect -1680 -35 -1672 -18
rect -2472 -59 -1672 -35
rect -1643 -18 -843 -10
rect -1643 -35 -1635 -18
rect -851 -35 -843 -18
rect -1643 -59 -843 -35
rect -814 -18 -14 -10
rect -814 -35 -806 -18
rect -22 -35 -14 -18
rect -814 -59 -14 -35
rect 14 -18 814 -10
rect 14 -35 22 -18
rect 806 -35 814 -18
rect 14 -59 814 -35
rect 843 -18 1643 -10
rect 843 -35 851 -18
rect 1635 -35 1643 -18
rect 843 -59 1643 -35
rect 1672 -18 2472 -10
rect 1672 -35 1680 -18
rect 2464 -35 2472 -18
rect 1672 -59 2472 -35
rect 2501 -18 3301 -10
rect 2501 -35 2509 -18
rect 3293 -35 3301 -18
rect 2501 -59 3301 -35
rect 3330 -18 4130 -10
rect 3330 -35 3338 -18
rect 4122 -35 4130 -18
rect 3330 -59 4130 -35
rect -4130 -124 -3330 -101
rect -4130 -141 -4122 -124
rect -3338 -141 -3330 -124
rect -4130 -149 -3330 -141
rect -3301 -124 -2501 -101
rect -3301 -141 -3293 -124
rect -2509 -141 -2501 -124
rect -3301 -149 -2501 -141
rect -2472 -124 -1672 -101
rect -2472 -141 -2464 -124
rect -1680 -141 -1672 -124
rect -2472 -149 -1672 -141
rect -1643 -124 -843 -101
rect -1643 -141 -1635 -124
rect -851 -141 -843 -124
rect -1643 -149 -843 -141
rect -814 -124 -14 -101
rect -814 -141 -806 -124
rect -22 -141 -14 -124
rect -814 -149 -14 -141
rect 14 -124 814 -101
rect 14 -141 22 -124
rect 806 -141 814 -124
rect 14 -149 814 -141
rect 843 -124 1643 -101
rect 843 -141 851 -124
rect 1635 -141 1643 -124
rect 843 -149 1643 -141
rect 1672 -124 2472 -101
rect 1672 -141 1680 -124
rect 2464 -141 2472 -124
rect 1672 -149 2472 -141
rect 2501 -124 3301 -101
rect 2501 -141 2509 -124
rect 3293 -141 3301 -124
rect 2501 -149 3301 -141
rect 3330 -124 4130 -101
rect 3330 -141 3338 -124
rect 4122 -141 4130 -124
rect 3330 -149 4130 -141
<< polycont >>
rect -4122 124 -3338 141
rect -3293 124 -2509 141
rect -2464 124 -1680 141
rect -1635 124 -851 141
rect -806 124 -22 141
rect 22 124 806 141
rect 851 124 1635 141
rect 1680 124 2464 141
rect 2509 124 3293 141
rect 3338 124 4122 141
rect -4122 18 -3338 35
rect -3293 18 -2509 35
rect -2464 18 -1680 35
rect -1635 18 -851 35
rect -806 18 -22 35
rect 22 18 806 35
rect 851 18 1635 35
rect 1680 18 2464 35
rect 2509 18 3293 35
rect 3338 18 4122 35
rect -4122 -35 -3338 -18
rect -3293 -35 -2509 -18
rect -2464 -35 -1680 -18
rect -1635 -35 -851 -18
rect -806 -35 -22 -18
rect 22 -35 806 -18
rect 851 -35 1635 -18
rect 1680 -35 2464 -18
rect 2509 -35 3293 -18
rect 3338 -35 4122 -18
rect -4122 -141 -3338 -124
rect -3293 -141 -2509 -124
rect -2464 -141 -1680 -124
rect -1635 -141 -851 -124
rect -806 -141 -22 -124
rect 22 -141 806 -124
rect 851 -141 1635 -124
rect 1680 -141 2464 -124
rect 2509 -141 3293 -124
rect 3338 -141 4122 -124
<< locali >>
rect -4220 193 -4172 210
rect 4172 193 4220 210
rect -4220 162 -4203 193
rect 4203 162 4220 193
rect -4130 124 -4122 141
rect -3338 124 -3330 141
rect -3301 124 -3293 141
rect -2509 124 -2501 141
rect -2472 124 -2464 141
rect -1680 124 -1672 141
rect -1643 124 -1635 141
rect -851 124 -843 141
rect -814 124 -806 141
rect -22 124 -14 141
rect 14 124 22 141
rect 806 124 814 141
rect 843 124 851 141
rect 1635 124 1643 141
rect 1672 124 1680 141
rect 2464 124 2472 141
rect 2501 124 2509 141
rect 3293 124 3301 141
rect 3330 124 3338 141
rect 4122 124 4130 141
rect -4153 95 -4136 103
rect -4153 57 -4136 65
rect -3324 95 -3307 103
rect -3324 57 -3307 65
rect -2495 95 -2478 103
rect -2495 57 -2478 65
rect -1666 95 -1649 103
rect -1666 57 -1649 65
rect -837 95 -820 103
rect -837 57 -820 65
rect -8 95 8 103
rect -8 57 8 65
rect 820 95 837 103
rect 820 57 837 65
rect 1649 95 1666 103
rect 1649 57 1666 65
rect 2478 95 2495 103
rect 2478 57 2495 65
rect 3307 95 3324 103
rect 3307 57 3324 65
rect 4136 95 4153 103
rect 4136 57 4153 65
rect -4130 18 -4122 35
rect -3338 18 -3330 35
rect -3301 18 -3293 35
rect -2509 18 -2501 35
rect -2472 18 -2464 35
rect -1680 18 -1672 35
rect -1643 18 -1635 35
rect -851 18 -843 35
rect -814 18 -806 35
rect -22 18 -14 35
rect 14 18 22 35
rect 806 18 814 35
rect 843 18 851 35
rect 1635 18 1643 35
rect 1672 18 1680 35
rect 2464 18 2472 35
rect 2501 18 2509 35
rect 3293 18 3301 35
rect 3330 18 3338 35
rect 4122 18 4130 35
rect -4130 -35 -4122 -18
rect -3338 -35 -3330 -18
rect -3301 -35 -3293 -18
rect -2509 -35 -2501 -18
rect -2472 -35 -2464 -18
rect -1680 -35 -1672 -18
rect -1643 -35 -1635 -18
rect -851 -35 -843 -18
rect -814 -35 -806 -18
rect -22 -35 -14 -18
rect 14 -35 22 -18
rect 806 -35 814 -18
rect 843 -35 851 -18
rect 1635 -35 1643 -18
rect 1672 -35 1680 -18
rect 2464 -35 2472 -18
rect 2501 -35 2509 -18
rect 3293 -35 3301 -18
rect 3330 -35 3338 -18
rect 4122 -35 4130 -18
rect -4153 -65 -4136 -57
rect -4153 -103 -4136 -95
rect -3324 -65 -3307 -57
rect -3324 -103 -3307 -95
rect -2495 -65 -2478 -57
rect -2495 -103 -2478 -95
rect -1666 -65 -1649 -57
rect -1666 -103 -1649 -95
rect -837 -65 -820 -57
rect -837 -103 -820 -95
rect -8 -65 8 -57
rect -8 -103 8 -95
rect 820 -65 837 -57
rect 820 -103 837 -95
rect 1649 -65 1666 -57
rect 1649 -103 1666 -95
rect 2478 -65 2495 -57
rect 2478 -103 2495 -95
rect 3307 -65 3324 -57
rect 3307 -103 3324 -95
rect 4136 -65 4153 -57
rect 4136 -103 4153 -95
rect -4130 -141 -4122 -124
rect -3338 -141 -3330 -124
rect -3301 -141 -3293 -124
rect -2509 -141 -2501 -124
rect -2472 -141 -2464 -124
rect -1680 -141 -1672 -124
rect -1643 -141 -1635 -124
rect -851 -141 -843 -124
rect -814 -141 -806 -124
rect -22 -141 -14 -124
rect 14 -141 22 -124
rect 806 -141 814 -124
rect 843 -141 851 -124
rect 1635 -141 1643 -124
rect 1672 -141 1680 -124
rect 2464 -141 2472 -124
rect 2501 -141 2509 -124
rect 3293 -141 3301 -124
rect 3330 -141 3338 -124
rect 4122 -141 4130 -124
rect -4220 -193 -4203 -162
rect 4203 -193 4220 -162
rect -4220 -210 -4172 -193
rect 4172 -210 4220 -193
<< viali >>
rect -4122 124 -3338 141
rect -3293 124 -2509 141
rect -2464 124 -1680 141
rect -1635 124 -851 141
rect -806 124 -22 141
rect 22 124 806 141
rect 851 124 1635 141
rect 1680 124 2464 141
rect 2509 124 3293 141
rect 3338 124 4122 141
rect -4153 65 -4136 95
rect -3324 65 -3307 95
rect -2495 65 -2478 95
rect -1666 65 -1649 95
rect -837 65 -820 95
rect -8 65 8 95
rect 820 65 837 95
rect 1649 65 1666 95
rect 2478 65 2495 95
rect 3307 65 3324 95
rect 4136 65 4153 95
rect -4122 18 -3338 35
rect -3293 18 -2509 35
rect -2464 18 -1680 35
rect -1635 18 -851 35
rect -806 18 -22 35
rect 22 18 806 35
rect 851 18 1635 35
rect 1680 18 2464 35
rect 2509 18 3293 35
rect 3338 18 4122 35
rect -4122 -35 -3338 -18
rect -3293 -35 -2509 -18
rect -2464 -35 -1680 -18
rect -1635 -35 -851 -18
rect -806 -35 -22 -18
rect 22 -35 806 -18
rect 851 -35 1635 -18
rect 1680 -35 2464 -18
rect 2509 -35 3293 -18
rect 3338 -35 4122 -18
rect -4153 -95 -4136 -65
rect -3324 -95 -3307 -65
rect -2495 -95 -2478 -65
rect -1666 -95 -1649 -65
rect -837 -95 -820 -65
rect -8 -95 8 -65
rect 820 -95 837 -65
rect 1649 -95 1666 -65
rect 2478 -95 2495 -65
rect 3307 -95 3324 -65
rect 4136 -95 4153 -65
rect -4122 -141 -3338 -124
rect -3293 -141 -2509 -124
rect -2464 -141 -1680 -124
rect -1635 -141 -851 -124
rect -806 -141 -22 -124
rect 22 -141 806 -124
rect 851 -141 1635 -124
rect 1680 -141 2464 -124
rect 2509 -141 3293 -124
rect 3338 -141 4122 -124
<< metal1 >>
rect -4128 141 -3332 144
rect -4128 124 -4122 141
rect -3338 124 -3332 141
rect -4128 121 -3332 124
rect -3299 141 -2503 144
rect -3299 124 -3293 141
rect -2509 124 -2503 141
rect -3299 121 -2503 124
rect -2470 141 -1674 144
rect -2470 124 -2464 141
rect -1680 124 -1674 141
rect -2470 121 -1674 124
rect -1641 141 -845 144
rect -1641 124 -1635 141
rect -851 124 -845 141
rect -1641 121 -845 124
rect -812 141 -16 144
rect -812 124 -806 141
rect -22 124 -16 141
rect -812 121 -16 124
rect 16 141 812 144
rect 16 124 22 141
rect 806 124 812 141
rect 16 121 812 124
rect 845 141 1641 144
rect 845 124 851 141
rect 1635 124 1641 141
rect 845 121 1641 124
rect 1674 141 2470 144
rect 1674 124 1680 141
rect 2464 124 2470 141
rect 1674 121 2470 124
rect 2503 141 3299 144
rect 2503 124 2509 141
rect 3293 124 3299 141
rect 2503 121 3299 124
rect 3332 141 4128 144
rect 3332 124 3338 141
rect 4122 124 4128 141
rect 3332 121 4128 124
rect -4156 95 -4133 101
rect -4156 65 -4153 95
rect -4136 65 -4133 95
rect -4156 59 -4133 65
rect -3327 95 -3304 101
rect -3327 65 -3324 95
rect -3307 65 -3304 95
rect -3327 59 -3304 65
rect -2498 95 -2475 101
rect -2498 65 -2495 95
rect -2478 65 -2475 95
rect -2498 59 -2475 65
rect -1669 95 -1646 101
rect -1669 65 -1666 95
rect -1649 65 -1646 95
rect -1669 59 -1646 65
rect -840 95 -817 101
rect -840 65 -837 95
rect -820 65 -817 95
rect -840 59 -817 65
rect -11 95 11 101
rect -11 65 -8 95
rect 8 65 11 95
rect -11 59 11 65
rect 817 95 840 101
rect 817 65 820 95
rect 837 65 840 95
rect 817 59 840 65
rect 1646 95 1669 101
rect 1646 65 1649 95
rect 1666 65 1669 95
rect 1646 59 1669 65
rect 2475 95 2498 101
rect 2475 65 2478 95
rect 2495 65 2498 95
rect 2475 59 2498 65
rect 3304 95 3327 101
rect 3304 65 3307 95
rect 3324 65 3327 95
rect 3304 59 3327 65
rect 4133 95 4156 101
rect 4133 65 4136 95
rect 4153 65 4156 95
rect 4133 59 4156 65
rect -4128 35 -3332 38
rect -4128 18 -4122 35
rect -3338 18 -3332 35
rect -4128 15 -3332 18
rect -3299 35 -2503 38
rect -3299 18 -3293 35
rect -2509 18 -2503 35
rect -3299 15 -2503 18
rect -2470 35 -1674 38
rect -2470 18 -2464 35
rect -1680 18 -1674 35
rect -2470 15 -1674 18
rect -1641 35 -845 38
rect -1641 18 -1635 35
rect -851 18 -845 35
rect -1641 15 -845 18
rect -812 35 -16 38
rect -812 18 -806 35
rect -22 18 -16 35
rect -812 15 -16 18
rect 16 35 812 38
rect 16 18 22 35
rect 806 18 812 35
rect 16 15 812 18
rect 845 35 1641 38
rect 845 18 851 35
rect 1635 18 1641 35
rect 845 15 1641 18
rect 1674 35 2470 38
rect 1674 18 1680 35
rect 2464 18 2470 35
rect 1674 15 2470 18
rect 2503 35 3299 38
rect 2503 18 2509 35
rect 3293 18 3299 35
rect 2503 15 3299 18
rect 3332 35 4128 38
rect 3332 18 3338 35
rect 4122 18 4128 35
rect 3332 15 4128 18
rect -4128 -18 -3332 -15
rect -4128 -35 -4122 -18
rect -3338 -35 -3332 -18
rect -4128 -38 -3332 -35
rect -3299 -18 -2503 -15
rect -3299 -35 -3293 -18
rect -2509 -35 -2503 -18
rect -3299 -38 -2503 -35
rect -2470 -18 -1674 -15
rect -2470 -35 -2464 -18
rect -1680 -35 -1674 -18
rect -2470 -38 -1674 -35
rect -1641 -18 -845 -15
rect -1641 -35 -1635 -18
rect -851 -35 -845 -18
rect -1641 -38 -845 -35
rect -812 -18 -16 -15
rect -812 -35 -806 -18
rect -22 -35 -16 -18
rect -812 -38 -16 -35
rect 16 -18 812 -15
rect 16 -35 22 -18
rect 806 -35 812 -18
rect 16 -38 812 -35
rect 845 -18 1641 -15
rect 845 -35 851 -18
rect 1635 -35 1641 -18
rect 845 -38 1641 -35
rect 1674 -18 2470 -15
rect 1674 -35 1680 -18
rect 2464 -35 2470 -18
rect 1674 -38 2470 -35
rect 2503 -18 3299 -15
rect 2503 -35 2509 -18
rect 3293 -35 3299 -18
rect 2503 -38 3299 -35
rect 3332 -18 4128 -15
rect 3332 -35 3338 -18
rect 4122 -35 4128 -18
rect 3332 -38 4128 -35
rect -4156 -65 -4133 -59
rect -4156 -95 -4153 -65
rect -4136 -95 -4133 -65
rect -4156 -101 -4133 -95
rect -3327 -65 -3304 -59
rect -3327 -95 -3324 -65
rect -3307 -95 -3304 -65
rect -3327 -101 -3304 -95
rect -2498 -65 -2475 -59
rect -2498 -95 -2495 -65
rect -2478 -95 -2475 -65
rect -2498 -101 -2475 -95
rect -1669 -65 -1646 -59
rect -1669 -95 -1666 -65
rect -1649 -95 -1646 -65
rect -1669 -101 -1646 -95
rect -840 -65 -817 -59
rect -840 -95 -837 -65
rect -820 -95 -817 -65
rect -840 -101 -817 -95
rect -11 -65 11 -59
rect -11 -95 -8 -65
rect 8 -95 11 -65
rect -11 -101 11 -95
rect 817 -65 840 -59
rect 817 -95 820 -65
rect 837 -95 840 -65
rect 817 -101 840 -95
rect 1646 -65 1669 -59
rect 1646 -95 1649 -65
rect 1666 -95 1669 -65
rect 1646 -101 1669 -95
rect 2475 -65 2498 -59
rect 2475 -95 2478 -65
rect 2495 -95 2498 -65
rect 2475 -101 2498 -95
rect 3304 -65 3327 -59
rect 3304 -95 3307 -65
rect 3324 -95 3327 -65
rect 3304 -101 3327 -95
rect 4133 -65 4156 -59
rect 4133 -95 4136 -65
rect 4153 -95 4156 -65
rect 4133 -101 4156 -95
rect -4128 -124 -3332 -121
rect -4128 -141 -4122 -124
rect -3338 -141 -3332 -124
rect -4128 -144 -3332 -141
rect -3299 -124 -2503 -121
rect -3299 -141 -3293 -124
rect -2509 -141 -2503 -124
rect -3299 -144 -2503 -141
rect -2470 -124 -1674 -121
rect -2470 -141 -2464 -124
rect -1680 -141 -1674 -124
rect -2470 -144 -1674 -141
rect -1641 -124 -845 -121
rect -1641 -141 -1635 -124
rect -851 -141 -845 -124
rect -1641 -144 -845 -141
rect -812 -124 -16 -121
rect -812 -141 -806 -124
rect -22 -141 -16 -124
rect -812 -144 -16 -141
rect 16 -124 812 -121
rect 16 -141 22 -124
rect 806 -141 812 -124
rect 16 -144 812 -141
rect 845 -124 1641 -121
rect 845 -141 851 -124
rect 1635 -141 1641 -124
rect 845 -144 1641 -141
rect 1674 -124 2470 -121
rect 1674 -141 1680 -124
rect 2464 -141 2470 -124
rect 1674 -144 2470 -141
rect 2503 -124 3299 -121
rect 2503 -141 2509 -124
rect 3293 -141 3299 -124
rect 2503 -144 3299 -141
rect 3332 -124 4128 -121
rect 3332 -141 3338 -124
rect 4122 -141 4128 -124
rect 3332 -144 4128 -141
<< properties >>
string FIXED_BBOX -4212 -202 4212 202
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 8.0 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
