magic
tech sky130A
magscale 1 2
timestamp 1712027638
<< pwell >>
rect -451 -4082 451 4082
<< psubdiff >>
rect -415 4012 -319 4046
rect 319 4012 415 4046
rect -415 3950 -381 4012
rect 381 3950 415 4012
rect -415 -4012 -381 -3950
rect 381 -4012 415 -3950
rect -415 -4046 -319 -4012
rect 319 -4046 415 -4012
<< psubdiffcont >>
rect -319 4012 319 4046
rect -415 -3950 -381 3950
rect 381 -3950 415 3950
rect -319 -4046 319 -4012
<< xpolycontact >>
rect -285 3484 285 3916
rect -285 -3916 285 -3484
<< xpolyres >>
rect -285 -3484 285 3484
<< locali >>
rect -415 4012 -319 4046
rect 319 4012 415 4046
rect -415 3950 -381 4012
rect 381 3950 415 4012
rect -415 -4012 -381 -3950
rect 381 -4012 415 -3950
rect -415 -4046 -319 -4012
rect 319 -4046 415 -4012
<< viali >>
rect -269 3501 269 3898
rect -269 -3898 269 -3501
<< metal1 >>
rect -281 3898 281 3904
rect -281 3501 -269 3898
rect 269 3501 281 3898
rect -281 3495 281 3501
rect -281 -3501 281 -3495
rect -281 -3898 -269 -3501
rect 269 -3898 281 -3501
rect -281 -3904 281 -3898
<< properties >>
string FIXED_BBOX -398 -4029 398 4029
string gencell sky130_fd_pr__res_xhigh_po_2p85
string library sky130
string parameters w 2.850 l 35 m 1 nx 1 wmin 2.850 lmin 0.50 rho 2000 val 24.693k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 2.850 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
