magic
tech sky130A
magscale 1 2
timestamp 1711677339
<< dnwell >>
rect 8363 -9837 36013 3064
<< nwell >>
rect 8283 2858 36093 3144
rect 8283 -9631 8569 2858
rect 35807 -9631 36093 2858
rect 8283 -9917 36093 -9631
<< pwell >>
rect 11372 -7488 31863 -896
<< nsubdiff >>
rect 8320 3087 36056 3107
rect 8320 3053 8400 3087
rect 35976 3053 36056 3087
rect 8320 3033 36056 3053
rect 8320 3027 8394 3033
rect 8320 -9800 8340 3027
rect 8374 -9800 8394 3027
rect 35982 3027 36056 3033
rect 8320 -9806 8394 -9800
rect 35982 -9800 36002 3027
rect 36036 -9800 36056 3027
rect 35982 -9806 36056 -9800
rect 8320 -9826 36056 -9806
rect 8320 -9860 8400 -9826
rect 35976 -9860 36056 -9826
rect 8320 -9880 36056 -9860
<< mvpsubdiff >>
rect 11952 -1660 31088 -1602
rect 11952 -2031 12010 -1660
rect 11952 -2081 11964 -2031
rect 11998 -2081 12010 -2031
rect 11952 -6681 12010 -2081
rect 31030 -6681 31088 -1660
rect 11952 -6739 31088 -6681
<< nsubdiffcont >>
rect 8400 3053 35976 3087
rect 8340 -9800 8374 3027
rect 36002 -9800 36036 3027
rect 8400 -9860 35976 -9826
<< mvpsubdiffcont >>
rect 11964 -2081 11998 -2031
<< locali >>
rect 8340 3053 8400 3087
rect 35976 3053 36036 3087
rect 8340 3027 8374 3053
rect 36002 3027 36036 3053
rect 11964 -1648 31076 -1614
rect 11964 -1892 11998 -1648
rect 11964 -2031 11998 -1957
rect 11964 -2255 11998 -2081
rect 11964 -3455 11998 -2289
rect 11964 -4655 11998 -3489
rect 11964 -5855 11998 -4689
rect 11964 -6727 11998 -5889
rect 8340 -9826 8374 -9800
rect 36002 -9826 36036 -9800
rect 8340 -9860 8400 -9826
rect 35976 -9860 36036 -9826
<< viali >>
rect 8340 -2485 8374 -2423
rect 11964 -1957 11998 -1892
rect 11964 -2289 11998 -2255
rect 11964 -3489 11998 -3455
rect 11964 -4689 11998 -4655
rect 11964 -5889 11998 -5855
<< metal1 >>
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 11953 -1892 12009 -1877
rect 11953 -1957 11964 -1892
rect 11998 -1957 12009 -1892
rect 18094 -1886 18150 -1880
rect 18094 -1948 18150 -1942
rect 19930 -1886 19986 -1880
rect 19930 -1948 19986 -1942
rect 23312 -1886 23368 -1880
rect 23312 -1948 23368 -1942
rect 25150 -1888 25202 -1882
rect 25150 -1946 25202 -1940
rect 11953 -2013 12009 -1957
rect 14422 -2004 14478 -1998
rect 14422 -2066 14478 -2060
rect 16258 -2004 16314 -1998
rect 16258 -2066 16314 -2060
rect 14256 -2119 14312 -2113
rect 14256 -2181 14312 -2175
rect 11952 -2255 12591 -2249
rect 11952 -2289 11964 -2255
rect 11998 -2289 12591 -2255
rect 11952 -2295 12591 -2289
rect 14183 -2295 14249 -2249
rect 14261 -2289 14307 -2181
rect 14427 -2295 14473 -2066
rect 16092 -2119 16148 -2113
rect 16092 -2181 16148 -2175
rect 16097 -2289 16143 -2181
rect 16263 -2295 16309 -2066
rect 17928 -2119 17984 -2113
rect 17928 -2181 17984 -2175
rect 17933 -2289 17979 -2181
rect 18099 -2295 18145 -1948
rect 19764 -2119 19820 -2113
rect 19764 -2181 19820 -2175
rect 19769 -2289 19815 -2181
rect 19935 -2295 19981 -1948
rect 21600 -2119 21656 -2113
rect 21600 -2181 21656 -2175
rect 21605 -2289 21651 -2181
rect 23317 -2295 23363 -1948
rect 23436 -2119 23492 -2113
rect 23436 -2181 23492 -2175
rect 23441 -2289 23487 -2181
rect 25153 -2295 25199 -1946
rect 26984 -2004 27040 -1998
rect 26984 -2066 27040 -2060
rect 28820 -2004 28876 -1998
rect 28820 -2066 28876 -2060
rect 25272 -2119 25328 -2113
rect 25272 -2181 25328 -2175
rect 25277 -2289 25323 -2181
rect 26989 -2295 27035 -2066
rect 27108 -2119 27164 -2113
rect 27108 -2181 27164 -2175
rect 27113 -2289 27159 -2181
rect 28825 -2295 28871 -2066
rect 28944 -2119 29000 -2113
rect 28944 -2181 29000 -2175
rect 28949 -2289 28995 -2181
rect 29049 -2295 29115 -2249
rect 30707 -2295 30763 -2249
rect 12535 -2327 12581 -2295
rect 30717 -2327 30763 -2295
rect 8329 -2423 8385 -2409
rect 8329 -2485 8340 -2423
rect 8374 -2485 8385 -2423
rect 8329 -2497 8385 -2485
rect 12535 -2494 12581 -2399
rect 14193 -2494 14239 -2399
rect 14371 -2494 14417 -2399
rect 12530 -2504 12586 -2494
rect 12530 -2570 12586 -2560
rect 14188 -2504 14244 -2494
rect 14188 -2570 14244 -2560
rect 14366 -2504 14422 -2494
rect 14366 -2570 14422 -2560
rect 16029 -2609 16075 -2411
rect 16207 -2494 16253 -2399
rect 16202 -2504 16258 -2494
rect 16202 -2570 16258 -2560
rect 17865 -2609 17911 -2411
rect 18043 -2494 18089 -2399
rect 18038 -2504 18094 -2494
rect 18038 -2570 18094 -2560
rect 16024 -2619 16080 -2609
rect 16024 -2685 16080 -2675
rect 17860 -2619 17916 -2609
rect 17860 -2685 17916 -2675
rect 19701 -2766 19747 -2411
rect 19879 -2494 19925 -2399
rect 19874 -2504 19930 -2494
rect 19874 -2570 19930 -2560
rect 21537 -2766 21583 -2399
rect 21715 -2766 21761 -2399
rect 23373 -2494 23419 -2399
rect 23368 -2504 23424 -2494
rect 23368 -2570 23424 -2560
rect 23551 -2766 23597 -2411
rect 25209 -2494 25255 -2399
rect 25204 -2504 25260 -2494
rect 25204 -2570 25260 -2560
rect 25387 -2609 25433 -2411
rect 27045 -2494 27091 -2399
rect 27040 -2504 27096 -2494
rect 27040 -2570 27096 -2560
rect 27223 -2609 27269 -2411
rect 28881 -2494 28927 -2399
rect 29059 -2494 29105 -2399
rect 30717 -2494 30763 -2399
rect 28876 -2504 28932 -2494
rect 28876 -2570 28932 -2560
rect 29054 -2504 29110 -2494
rect 29054 -2570 29110 -2560
rect 30712 -2504 30768 -2494
rect 30712 -2570 30768 -2560
rect 25382 -2619 25438 -2609
rect 25382 -2685 25438 -2675
rect 27218 -2619 27274 -2609
rect 27218 -2685 27274 -2675
rect 19686 -2822 19696 -2766
rect 19752 -2822 19762 -2766
rect 21522 -2822 21532 -2766
rect 21588 -2822 21598 -2766
rect 21700 -2822 21710 -2766
rect 21766 -2822 21776 -2766
rect 23536 -2822 23546 -2766
rect 23602 -2822 23612 -2766
rect 18094 -3086 18150 -3080
rect 18094 -3148 18150 -3142
rect 19930 -3086 19986 -3080
rect 19930 -3148 19986 -3142
rect 23312 -3086 23368 -3080
rect 23312 -3148 23368 -3142
rect 25150 -3088 25202 -3082
rect 25150 -3146 25202 -3140
rect 14422 -3204 14478 -3198
rect 14422 -3266 14478 -3260
rect 16258 -3204 16314 -3198
rect 16258 -3266 16314 -3260
rect 14256 -3319 14312 -3313
rect 14256 -3381 14312 -3375
rect 11952 -3455 12591 -3449
rect 11952 -3489 11964 -3455
rect 11998 -3489 12591 -3455
rect 11952 -3495 12591 -3489
rect 14183 -3495 14249 -3449
rect 14261 -3489 14307 -3381
rect 14427 -3495 14473 -3266
rect 16092 -3319 16148 -3313
rect 16092 -3381 16148 -3375
rect 16097 -3489 16143 -3381
rect 16263 -3495 16309 -3266
rect 17928 -3319 17984 -3313
rect 17928 -3381 17984 -3375
rect 17933 -3489 17979 -3381
rect 18099 -3495 18145 -3148
rect 19764 -3319 19820 -3313
rect 19764 -3381 19820 -3375
rect 19769 -3489 19815 -3381
rect 19935 -3495 19981 -3148
rect 21600 -3319 21656 -3313
rect 21600 -3381 21656 -3375
rect 21605 -3489 21651 -3381
rect 23317 -3495 23363 -3148
rect 23436 -3319 23492 -3313
rect 23436 -3381 23492 -3375
rect 23441 -3489 23487 -3381
rect 25153 -3495 25199 -3146
rect 26984 -3204 27040 -3198
rect 26984 -3266 27040 -3260
rect 28820 -3204 28876 -3198
rect 28820 -3266 28876 -3260
rect 25272 -3319 25328 -3313
rect 25272 -3381 25328 -3375
rect 25277 -3489 25323 -3381
rect 26989 -3495 27035 -3266
rect 27108 -3319 27164 -3313
rect 27108 -3381 27164 -3375
rect 27113 -3489 27159 -3381
rect 28825 -3495 28871 -3266
rect 28944 -3319 29000 -3313
rect 28944 -3381 29000 -3375
rect 28949 -3489 28995 -3381
rect 29049 -3495 29115 -3449
rect 30707 -3495 30763 -3449
rect 12535 -3527 12581 -3495
rect 30717 -3527 30763 -3495
rect 12535 -3694 12581 -3599
rect 14193 -3694 14239 -3599
rect 14371 -3694 14417 -3599
rect 12530 -3704 12586 -3694
rect 12530 -3770 12586 -3760
rect 14188 -3704 14244 -3694
rect 14188 -3770 14244 -3760
rect 14366 -3704 14422 -3694
rect 14366 -3770 14422 -3760
rect 16029 -3809 16075 -3611
rect 16207 -3694 16253 -3599
rect 16202 -3704 16258 -3694
rect 16202 -3770 16258 -3760
rect 17865 -3809 17911 -3611
rect 18043 -3694 18089 -3599
rect 18038 -3704 18094 -3694
rect 18038 -3770 18094 -3760
rect 16024 -3819 16080 -3809
rect 16024 -3885 16080 -3875
rect 17860 -3819 17916 -3809
rect 17860 -3885 17916 -3875
rect 19701 -3966 19747 -3611
rect 19879 -3694 19925 -3599
rect 19874 -3704 19930 -3694
rect 19874 -3770 19930 -3760
rect 21537 -3966 21583 -3599
rect 21715 -3966 21761 -3599
rect 23373 -3694 23419 -3599
rect 23368 -3704 23424 -3694
rect 23368 -3770 23424 -3760
rect 23551 -3966 23597 -3611
rect 25209 -3694 25255 -3599
rect 25204 -3704 25260 -3694
rect 25204 -3770 25260 -3760
rect 25387 -3809 25433 -3611
rect 27045 -3694 27091 -3599
rect 27040 -3704 27096 -3694
rect 27040 -3770 27096 -3760
rect 27223 -3809 27269 -3611
rect 28881 -3694 28927 -3599
rect 29059 -3694 29105 -3599
rect 30717 -3694 30763 -3599
rect 28876 -3704 28932 -3694
rect 28876 -3770 28932 -3760
rect 29054 -3704 29110 -3694
rect 29054 -3770 29110 -3760
rect 30712 -3704 30768 -3694
rect 30712 -3770 30768 -3760
rect 25382 -3819 25438 -3809
rect 25382 -3885 25438 -3875
rect 27218 -3819 27274 -3809
rect 27218 -3885 27274 -3875
rect 19686 -4022 19696 -3966
rect 19752 -4022 19762 -3966
rect 21522 -4022 21532 -3966
rect 21588 -4022 21598 -3966
rect 21700 -4022 21710 -3966
rect 21766 -4022 21776 -3966
rect 23536 -4022 23546 -3966
rect 23602 -4022 23612 -3966
rect 18094 -4286 18150 -4280
rect 18094 -4348 18150 -4342
rect 19930 -4286 19986 -4280
rect 19930 -4348 19986 -4342
rect 23312 -4286 23368 -4280
rect 23312 -4348 23368 -4342
rect 25150 -4288 25202 -4282
rect 25150 -4346 25202 -4340
rect 14422 -4404 14478 -4398
rect 14422 -4466 14478 -4460
rect 16258 -4404 16314 -4398
rect 16258 -4466 16314 -4460
rect 14256 -4519 14312 -4513
rect 14256 -4581 14312 -4575
rect 11952 -4655 12591 -4649
rect 11952 -4689 11964 -4655
rect 11998 -4689 12591 -4655
rect 11952 -4695 12591 -4689
rect 14183 -4695 14249 -4649
rect 14261 -4689 14307 -4581
rect 14427 -4695 14473 -4466
rect 16092 -4519 16148 -4513
rect 16092 -4581 16148 -4575
rect 16097 -4689 16143 -4581
rect 16263 -4695 16309 -4466
rect 17928 -4519 17984 -4513
rect 17928 -4581 17984 -4575
rect 17933 -4689 17979 -4581
rect 18099 -4695 18145 -4348
rect 19764 -4519 19820 -4513
rect 19764 -4581 19820 -4575
rect 19769 -4689 19815 -4581
rect 19935 -4695 19981 -4348
rect 21600 -4519 21656 -4513
rect 21600 -4581 21656 -4575
rect 21605 -4689 21651 -4581
rect 23317 -4695 23363 -4348
rect 23436 -4519 23492 -4513
rect 23436 -4581 23492 -4575
rect 23441 -4689 23487 -4581
rect 25153 -4695 25199 -4346
rect 26984 -4404 27040 -4398
rect 26984 -4466 27040 -4460
rect 28820 -4404 28876 -4398
rect 28820 -4466 28876 -4460
rect 25272 -4519 25328 -4513
rect 25272 -4581 25328 -4575
rect 25277 -4689 25323 -4581
rect 26989 -4695 27035 -4466
rect 27108 -4519 27164 -4513
rect 27108 -4581 27164 -4575
rect 27113 -4689 27159 -4581
rect 28825 -4695 28871 -4466
rect 28944 -4519 29000 -4513
rect 28944 -4581 29000 -4575
rect 28949 -4689 28995 -4581
rect 29049 -4695 29115 -4649
rect 30707 -4695 30763 -4649
rect 12535 -4727 12581 -4695
rect 30717 -4727 30763 -4695
rect 12535 -4894 12581 -4799
rect 14193 -4894 14239 -4799
rect 14371 -4894 14417 -4799
rect 12530 -4904 12586 -4894
rect 12530 -4970 12586 -4960
rect 14188 -4904 14244 -4894
rect 14188 -4970 14244 -4960
rect 14366 -4904 14422 -4894
rect 14366 -4970 14422 -4960
rect 16029 -5009 16075 -4811
rect 16207 -4894 16253 -4799
rect 16202 -4904 16258 -4894
rect 16202 -4970 16258 -4960
rect 17865 -5009 17911 -4811
rect 18043 -4894 18089 -4799
rect 18038 -4904 18094 -4894
rect 18038 -4970 18094 -4960
rect 16024 -5019 16080 -5009
rect 16024 -5085 16080 -5075
rect 17860 -5019 17916 -5009
rect 17860 -5085 17916 -5075
rect 19701 -5166 19747 -4811
rect 19879 -4894 19925 -4799
rect 19874 -4904 19930 -4894
rect 19874 -4970 19930 -4960
rect 21537 -5166 21583 -4799
rect 21715 -5166 21761 -4799
rect 23373 -4894 23419 -4799
rect 23368 -4904 23424 -4894
rect 23368 -4970 23424 -4960
rect 23551 -5166 23597 -4811
rect 25209 -4894 25255 -4799
rect 25204 -4904 25260 -4894
rect 25204 -4970 25260 -4960
rect 25387 -5009 25433 -4811
rect 27045 -4894 27091 -4799
rect 27040 -4904 27096 -4894
rect 27040 -4970 27096 -4960
rect 27223 -5009 27269 -4811
rect 28881 -4894 28927 -4799
rect 29059 -4894 29105 -4799
rect 30717 -4894 30763 -4799
rect 28876 -4904 28932 -4894
rect 28876 -4970 28932 -4960
rect 29054 -4904 29110 -4894
rect 29054 -4970 29110 -4960
rect 30712 -4904 30768 -4894
rect 30712 -4970 30768 -4960
rect 25382 -5019 25438 -5009
rect 25382 -5085 25438 -5075
rect 27218 -5019 27274 -5009
rect 27218 -5085 27274 -5075
rect 19686 -5222 19696 -5166
rect 19752 -5222 19762 -5166
rect 21522 -5222 21532 -5166
rect 21588 -5222 21598 -5166
rect 21700 -5222 21710 -5166
rect 21766 -5222 21776 -5166
rect 23536 -5222 23546 -5166
rect 23602 -5222 23612 -5166
rect 18094 -5486 18150 -5480
rect 18094 -5548 18150 -5542
rect 19930 -5486 19986 -5480
rect 19930 -5548 19986 -5542
rect 23312 -5486 23368 -5480
rect 23312 -5548 23368 -5542
rect 25150 -5488 25202 -5482
rect 25150 -5546 25202 -5540
rect 14422 -5604 14478 -5598
rect 14422 -5666 14478 -5660
rect 16258 -5604 16314 -5598
rect 16258 -5666 16314 -5660
rect 14256 -5719 14312 -5713
rect 14256 -5781 14312 -5775
rect 11952 -5855 12591 -5849
rect 11952 -5889 11964 -5855
rect 11998 -5889 12591 -5855
rect 11952 -5895 12591 -5889
rect 14183 -5895 14249 -5849
rect 14261 -5889 14307 -5781
rect 14427 -5895 14473 -5666
rect 16092 -5719 16148 -5713
rect 16092 -5781 16148 -5775
rect 16097 -5889 16143 -5781
rect 16263 -5895 16309 -5666
rect 17928 -5719 17984 -5713
rect 17928 -5781 17984 -5775
rect 17933 -5889 17979 -5781
rect 18099 -5895 18145 -5548
rect 19764 -5719 19820 -5713
rect 19764 -5781 19820 -5775
rect 19769 -5889 19815 -5781
rect 19935 -5895 19981 -5548
rect 21600 -5719 21656 -5713
rect 21600 -5781 21656 -5775
rect 21605 -5889 21651 -5781
rect 23317 -5895 23363 -5548
rect 23436 -5719 23492 -5713
rect 23436 -5781 23492 -5775
rect 23441 -5889 23487 -5781
rect 25153 -5895 25199 -5546
rect 26984 -5604 27040 -5598
rect 26984 -5666 27040 -5660
rect 28820 -5604 28876 -5598
rect 28820 -5666 28876 -5660
rect 25272 -5719 25328 -5713
rect 25272 -5781 25328 -5775
rect 25277 -5889 25323 -5781
rect 26989 -5895 27035 -5666
rect 27108 -5719 27164 -5713
rect 27108 -5781 27164 -5775
rect 27113 -5889 27159 -5781
rect 28825 -5895 28871 -5666
rect 28944 -5719 29000 -5713
rect 28944 -5781 29000 -5775
rect 28949 -5889 28995 -5781
rect 29049 -5895 29115 -5849
rect 30707 -5895 30763 -5849
rect 12535 -5927 12581 -5895
rect 30717 -5927 30763 -5895
rect 12535 -6094 12581 -5999
rect 14193 -6094 14239 -5999
rect 14371 -6094 14417 -5999
rect 12530 -6104 12586 -6094
rect 12530 -6170 12586 -6160
rect 14188 -6104 14244 -6094
rect 14188 -6170 14244 -6160
rect 14366 -6104 14422 -6094
rect 14366 -6170 14422 -6160
rect 16029 -6209 16075 -6011
rect 16207 -6094 16253 -5999
rect 16202 -6104 16258 -6094
rect 16202 -6170 16258 -6160
rect 17865 -6209 17911 -6011
rect 18043 -6094 18089 -5999
rect 18038 -6104 18094 -6094
rect 18038 -6170 18094 -6160
rect 16024 -6219 16080 -6209
rect 16024 -6285 16080 -6275
rect 17860 -6219 17916 -6209
rect 17860 -6285 17916 -6275
rect 19701 -6366 19747 -6011
rect 19879 -6094 19925 -5999
rect 19874 -6104 19930 -6094
rect 19874 -6170 19930 -6160
rect 21537 -6366 21583 -5999
rect 21715 -6366 21761 -5999
rect 23373 -6094 23419 -5999
rect 23368 -6104 23424 -6094
rect 23368 -6170 23424 -6160
rect 23551 -6366 23597 -6011
rect 25209 -6094 25255 -5999
rect 25204 -6104 25260 -6094
rect 25204 -6170 25260 -6160
rect 25387 -6209 25433 -6011
rect 27045 -6094 27091 -5999
rect 27040 -6104 27096 -6094
rect 27040 -6170 27096 -6160
rect 27223 -6209 27269 -6011
rect 28881 -6094 28927 -5999
rect 29059 -6094 29105 -5999
rect 30717 -6094 30763 -5999
rect 28876 -6104 28932 -6094
rect 28876 -6170 28932 -6160
rect 29054 -6104 29110 -6094
rect 29054 -6170 29110 -6160
rect 30712 -6104 30768 -6094
rect 30712 -6170 30768 -6160
rect 25382 -6219 25438 -6209
rect 25382 -6285 25438 -6275
rect 27218 -6219 27274 -6209
rect 27218 -6285 27274 -6275
rect 19686 -6422 19696 -6366
rect 19752 -6422 19762 -6366
rect 21522 -6422 21532 -6366
rect 21588 -6422 21598 -6366
rect 21700 -6422 21710 -6366
rect 21766 -6422 21776 -6366
rect 23536 -6422 23546 -6366
rect 23602 -6422 23612 -6366
<< via1 >>
rect 18094 -1942 18150 -1886
rect 19930 -1942 19986 -1886
rect 23312 -1942 23368 -1886
rect 25150 -1940 25202 -1888
rect 14422 -2060 14478 -2004
rect 16258 -2060 16314 -2004
rect 14256 -2175 14312 -2119
rect 16092 -2175 16148 -2119
rect 17928 -2175 17984 -2119
rect 19764 -2175 19820 -2119
rect 21600 -2175 21656 -2119
rect 23436 -2175 23492 -2119
rect 26984 -2060 27040 -2004
rect 28820 -2060 28876 -2004
rect 25272 -2175 25328 -2119
rect 27108 -2175 27164 -2119
rect 28944 -2175 29000 -2119
rect 12530 -2560 12586 -2504
rect 14188 -2560 14244 -2504
rect 14366 -2560 14422 -2504
rect 16202 -2560 16258 -2504
rect 18038 -2560 18094 -2504
rect 16024 -2675 16080 -2619
rect 17860 -2675 17916 -2619
rect 19874 -2560 19930 -2504
rect 23368 -2560 23424 -2504
rect 25204 -2560 25260 -2504
rect 27040 -2560 27096 -2504
rect 28876 -2560 28932 -2504
rect 29054 -2560 29110 -2504
rect 30712 -2560 30768 -2504
rect 25382 -2675 25438 -2619
rect 27218 -2675 27274 -2619
rect 19696 -2822 19752 -2766
rect 21532 -2822 21588 -2766
rect 21710 -2822 21766 -2766
rect 23546 -2822 23602 -2766
rect 18094 -3142 18150 -3086
rect 19930 -3142 19986 -3086
rect 23312 -3142 23368 -3086
rect 25150 -3140 25202 -3088
rect 14422 -3260 14478 -3204
rect 16258 -3260 16314 -3204
rect 14256 -3375 14312 -3319
rect 16092 -3375 16148 -3319
rect 17928 -3375 17984 -3319
rect 19764 -3375 19820 -3319
rect 21600 -3375 21656 -3319
rect 23436 -3375 23492 -3319
rect 26984 -3260 27040 -3204
rect 28820 -3260 28876 -3204
rect 25272 -3375 25328 -3319
rect 27108 -3375 27164 -3319
rect 28944 -3375 29000 -3319
rect 12530 -3760 12586 -3704
rect 14188 -3760 14244 -3704
rect 14366 -3760 14422 -3704
rect 16202 -3760 16258 -3704
rect 18038 -3760 18094 -3704
rect 16024 -3875 16080 -3819
rect 17860 -3875 17916 -3819
rect 19874 -3760 19930 -3704
rect 23368 -3760 23424 -3704
rect 25204 -3760 25260 -3704
rect 27040 -3760 27096 -3704
rect 28876 -3760 28932 -3704
rect 29054 -3760 29110 -3704
rect 30712 -3760 30768 -3704
rect 25382 -3875 25438 -3819
rect 27218 -3875 27274 -3819
rect 19696 -4022 19752 -3966
rect 21532 -4022 21588 -3966
rect 21710 -4022 21766 -3966
rect 23546 -4022 23602 -3966
rect 18094 -4342 18150 -4286
rect 19930 -4342 19986 -4286
rect 23312 -4342 23368 -4286
rect 25150 -4340 25202 -4288
rect 14422 -4460 14478 -4404
rect 16258 -4460 16314 -4404
rect 14256 -4575 14312 -4519
rect 16092 -4575 16148 -4519
rect 17928 -4575 17984 -4519
rect 19764 -4575 19820 -4519
rect 21600 -4575 21656 -4519
rect 23436 -4575 23492 -4519
rect 26984 -4460 27040 -4404
rect 28820 -4460 28876 -4404
rect 25272 -4575 25328 -4519
rect 27108 -4575 27164 -4519
rect 28944 -4575 29000 -4519
rect 12530 -4960 12586 -4904
rect 14188 -4960 14244 -4904
rect 14366 -4960 14422 -4904
rect 16202 -4960 16258 -4904
rect 18038 -4960 18094 -4904
rect 16024 -5075 16080 -5019
rect 17860 -5075 17916 -5019
rect 19874 -4960 19930 -4904
rect 23368 -4960 23424 -4904
rect 25204 -4960 25260 -4904
rect 27040 -4960 27096 -4904
rect 28876 -4960 28932 -4904
rect 29054 -4960 29110 -4904
rect 30712 -4960 30768 -4904
rect 25382 -5075 25438 -5019
rect 27218 -5075 27274 -5019
rect 19696 -5222 19752 -5166
rect 21532 -5222 21588 -5166
rect 21710 -5222 21766 -5166
rect 23546 -5222 23602 -5166
rect 18094 -5542 18150 -5486
rect 19930 -5542 19986 -5486
rect 23312 -5542 23368 -5486
rect 25150 -5540 25202 -5488
rect 14422 -5660 14478 -5604
rect 16258 -5660 16314 -5604
rect 14256 -5775 14312 -5719
rect 16092 -5775 16148 -5719
rect 17928 -5775 17984 -5719
rect 19764 -5775 19820 -5719
rect 21600 -5775 21656 -5719
rect 23436 -5775 23492 -5719
rect 26984 -5660 27040 -5604
rect 28820 -5660 28876 -5604
rect 25272 -5775 25328 -5719
rect 27108 -5775 27164 -5719
rect 28944 -5775 29000 -5719
rect 12530 -6160 12586 -6104
rect 14188 -6160 14244 -6104
rect 14366 -6160 14422 -6104
rect 16202 -6160 16258 -6104
rect 18038 -6160 18094 -6104
rect 16024 -6275 16080 -6219
rect 17860 -6275 17916 -6219
rect 19874 -6160 19930 -6104
rect 23368 -6160 23424 -6104
rect 25204 -6160 25260 -6104
rect 27040 -6160 27096 -6104
rect 28876 -6160 28932 -6104
rect 29054 -6160 29110 -6104
rect 30712 -6160 30768 -6104
rect 25382 -6275 25438 -6219
rect 27218 -6275 27274 -6219
rect 19696 -6422 19752 -6366
rect 21532 -6422 21588 -6366
rect 21710 -6422 21766 -6366
rect 23546 -6422 23602 -6366
<< metal2 >>
rect 18088 -1942 18094 -1886
rect 18150 -1942 19930 -1886
rect 19986 -1942 22482 -1886
rect 22538 -1942 23312 -1886
rect 23368 -1888 25208 -1886
rect 23368 -1940 25150 -1888
rect 25202 -1940 25208 -1888
rect 23368 -1942 25208 -1940
rect 14416 -2060 14422 -2004
rect 14478 -2060 16258 -2004
rect 16314 -2060 22266 -2004
rect 22322 -2060 26984 -2004
rect 27040 -2060 28820 -2004
rect 28876 -2060 28882 -2004
rect 14250 -2175 14256 -2119
rect 14312 -2175 16092 -2119
rect 16148 -2175 17928 -2119
rect 17984 -2175 19764 -2119
rect 19820 -2175 21600 -2119
rect 21656 -2175 23436 -2119
rect 23492 -2175 25272 -2119
rect 25328 -2175 27108 -2119
rect 27164 -2175 28944 -2119
rect 29000 -2175 29006 -2119
rect 12520 -2560 12530 -2504
rect 12586 -2560 14188 -2504
rect 14244 -2560 14254 -2504
rect 14360 -2560 14366 -2504
rect 14422 -2560 16202 -2504
rect 16258 -2560 18038 -2504
rect 18094 -2560 19874 -2504
rect 19930 -2560 20487 -2504
rect 20543 -2560 23368 -2504
rect 23424 -2560 25204 -2504
rect 25260 -2560 27040 -2504
rect 27096 -2560 28876 -2504
rect 28932 -2560 28942 -2504
rect 29044 -2560 29054 -2504
rect 29110 -2560 30712 -2504
rect 30768 -2560 30778 -2504
rect 16018 -2675 16024 -2619
rect 16080 -2675 17860 -2619
rect 17916 -2675 21147 -2619
rect 21203 -2675 25382 -2619
rect 25438 -2675 27218 -2619
rect 27274 -2675 27284 -2619
rect 19696 -2766 19752 -2756
rect 21532 -2766 21588 -2756
rect 21710 -2766 21766 -2756
rect 23546 -2766 23602 -2756
rect 19752 -2822 21346 -2766
rect 21402 -2822 21532 -2766
rect 21588 -2822 21710 -2766
rect 21766 -2822 23546 -2766
rect 19696 -2832 19752 -2822
rect 21532 -2832 21588 -2822
rect 21710 -2832 21766 -2822
rect 23546 -2832 23602 -2822
rect 18088 -3142 18094 -3086
rect 18150 -3142 19930 -3086
rect 19986 -3142 22482 -3086
rect 22538 -3142 23312 -3086
rect 23368 -3088 25208 -3086
rect 23368 -3140 25150 -3088
rect 25202 -3140 25208 -3088
rect 23368 -3142 25208 -3140
rect 14416 -3260 14422 -3204
rect 14478 -3260 16258 -3204
rect 16314 -3260 22266 -3204
rect 22322 -3260 26984 -3204
rect 27040 -3260 28820 -3204
rect 28876 -3260 28882 -3204
rect 14250 -3375 14256 -3319
rect 14312 -3375 16092 -3319
rect 16148 -3375 17928 -3319
rect 17984 -3375 19764 -3319
rect 19820 -3375 21600 -3319
rect 21656 -3375 23436 -3319
rect 23492 -3375 25272 -3319
rect 25328 -3375 27108 -3319
rect 27164 -3375 28944 -3319
rect 29000 -3375 29006 -3319
rect 12520 -3760 12530 -3704
rect 12586 -3760 14188 -3704
rect 14244 -3760 14254 -3704
rect 14360 -3760 14366 -3704
rect 14422 -3760 16202 -3704
rect 16258 -3760 18038 -3704
rect 18094 -3760 19874 -3704
rect 19930 -3760 20487 -3704
rect 20543 -3760 23368 -3704
rect 23424 -3760 25204 -3704
rect 25260 -3760 27040 -3704
rect 27096 -3760 28876 -3704
rect 28932 -3760 28942 -3704
rect 29044 -3760 29054 -3704
rect 29110 -3760 30712 -3704
rect 30768 -3760 30778 -3704
rect 16018 -3875 16024 -3819
rect 16080 -3875 17860 -3819
rect 17916 -3875 21147 -3819
rect 21203 -3875 25382 -3819
rect 25438 -3875 27218 -3819
rect 27274 -3875 27284 -3819
rect 19696 -3966 19752 -3956
rect 21532 -3966 21588 -3956
rect 21710 -3966 21766 -3956
rect 23546 -3966 23602 -3956
rect 19752 -4022 21346 -3966
rect 21402 -4022 21532 -3966
rect 21588 -4022 21710 -3966
rect 21766 -4022 23546 -3966
rect 19696 -4032 19752 -4022
rect 21532 -4032 21588 -4022
rect 21710 -4032 21766 -4022
rect 23546 -4032 23602 -4022
rect 18088 -4342 18094 -4286
rect 18150 -4342 19930 -4286
rect 19986 -4342 22482 -4286
rect 22538 -4342 23312 -4286
rect 23368 -4288 25208 -4286
rect 23368 -4340 25150 -4288
rect 25202 -4340 25208 -4288
rect 23368 -4342 25208 -4340
rect 14416 -4460 14422 -4404
rect 14478 -4460 16258 -4404
rect 16314 -4460 22266 -4404
rect 22322 -4460 26984 -4404
rect 27040 -4460 28820 -4404
rect 28876 -4460 28882 -4404
rect 14250 -4575 14256 -4519
rect 14312 -4575 16092 -4519
rect 16148 -4575 17928 -4519
rect 17984 -4575 19764 -4519
rect 19820 -4575 21600 -4519
rect 21656 -4575 23436 -4519
rect 23492 -4575 25272 -4519
rect 25328 -4575 27108 -4519
rect 27164 -4575 28944 -4519
rect 29000 -4575 29006 -4519
rect 12520 -4960 12530 -4904
rect 12586 -4960 14188 -4904
rect 14244 -4960 14254 -4904
rect 14360 -4960 14366 -4904
rect 14422 -4960 16202 -4904
rect 16258 -4960 18038 -4904
rect 18094 -4960 19874 -4904
rect 19930 -4960 20487 -4904
rect 20543 -4960 23368 -4904
rect 23424 -4960 25204 -4904
rect 25260 -4960 27040 -4904
rect 27096 -4960 28876 -4904
rect 28932 -4960 28942 -4904
rect 29044 -4960 29054 -4904
rect 29110 -4960 30712 -4904
rect 30768 -4960 30778 -4904
rect 16018 -5075 16024 -5019
rect 16080 -5075 17860 -5019
rect 17916 -5075 21147 -5019
rect 21203 -5075 25382 -5019
rect 25438 -5075 27218 -5019
rect 27274 -5075 27284 -5019
rect 19696 -5166 19752 -5156
rect 21532 -5166 21588 -5156
rect 21710 -5166 21766 -5156
rect 23546 -5166 23602 -5156
rect 19752 -5222 21346 -5166
rect 21402 -5222 21532 -5166
rect 21588 -5222 21710 -5166
rect 21766 -5222 23546 -5166
rect 19696 -5232 19752 -5222
rect 21532 -5232 21588 -5222
rect 21710 -5232 21766 -5222
rect 23546 -5232 23602 -5222
rect 18088 -5542 18094 -5486
rect 18150 -5542 19930 -5486
rect 19986 -5542 22482 -5486
rect 22538 -5542 23312 -5486
rect 23368 -5488 25208 -5486
rect 23368 -5540 25150 -5488
rect 25202 -5540 25208 -5488
rect 23368 -5542 25208 -5540
rect 14416 -5660 14422 -5604
rect 14478 -5660 16258 -5604
rect 16314 -5660 22266 -5604
rect 22322 -5660 26984 -5604
rect 27040 -5660 28820 -5604
rect 28876 -5660 28882 -5604
rect 14250 -5775 14256 -5719
rect 14312 -5775 16092 -5719
rect 16148 -5775 17928 -5719
rect 17984 -5775 19764 -5719
rect 19820 -5775 21600 -5719
rect 21656 -5775 23436 -5719
rect 23492 -5775 25272 -5719
rect 25328 -5775 27108 -5719
rect 27164 -5775 28944 -5719
rect 29000 -5775 29006 -5719
rect 12520 -6160 12530 -6104
rect 12586 -6160 14188 -6104
rect 14244 -6160 14254 -6104
rect 14360 -6160 14366 -6104
rect 14422 -6160 16202 -6104
rect 16258 -6160 18038 -6104
rect 18094 -6160 19874 -6104
rect 19930 -6160 20487 -6104
rect 20543 -6160 23368 -6104
rect 23424 -6160 25204 -6104
rect 25260 -6160 27040 -6104
rect 27096 -6160 28876 -6104
rect 28932 -6160 28942 -6104
rect 29044 -6160 29054 -6104
rect 29110 -6160 30712 -6104
rect 30768 -6160 30778 -6104
rect 16018 -6275 16024 -6219
rect 16080 -6275 17860 -6219
rect 17916 -6275 21147 -6219
rect 21203 -6275 25382 -6219
rect 25438 -6275 27218 -6219
rect 27274 -6275 27284 -6219
rect 19696 -6366 19752 -6356
rect 21532 -6366 21588 -6356
rect 21710 -6366 21766 -6356
rect 23546 -6366 23602 -6356
rect 19752 -6422 21346 -6366
rect 21402 -6422 21532 -6366
rect 21588 -6422 21710 -6366
rect 21766 -6422 23546 -6366
rect 19696 -6432 19752 -6422
rect 21532 -6432 21588 -6422
rect 21710 -6432 21766 -6422
rect 23546 -6432 23602 -6422
<< via2 >>
rect 22482 -1942 22538 -1886
rect 22266 -2060 22322 -2004
rect 20487 -2560 20543 -2504
rect 21147 -2675 21203 -2619
rect 21346 -2822 21402 -2766
rect 22482 -3142 22538 -3086
rect 22266 -3260 22322 -3204
rect 20487 -3760 20543 -3704
rect 21147 -3875 21203 -3819
rect 21346 -4022 21402 -3966
rect 22482 -4342 22538 -4286
rect 22266 -4460 22322 -4404
rect 20487 -4960 20543 -4904
rect 21147 -5075 21203 -5019
rect 21346 -5222 21402 -5166
rect 22482 -5542 22538 -5486
rect 22266 -5660 22322 -5604
rect 20487 -6160 20543 -6104
rect 21147 -6275 21203 -6219
rect 21346 -6422 21402 -6366
<< metal3 >>
rect 22472 -1886 22548 -1881
rect 22472 -1942 22482 -1886
rect 22538 -1942 22548 -1886
rect 22256 -2004 22332 -1999
rect 22256 -2060 22266 -2004
rect 22322 -2060 22332 -2004
rect 20477 -2504 20553 -2499
rect 20477 -2560 20487 -2504
rect 20543 -2560 20553 -2504
rect 20477 -3704 20553 -2560
rect 20477 -3760 20487 -3704
rect 20543 -3760 20553 -3704
rect 20477 -4904 20553 -3760
rect 20477 -4960 20487 -4904
rect 20543 -4960 20553 -4904
rect 20477 -6104 20553 -4960
rect 20477 -6160 20487 -6104
rect 20543 -6160 20553 -6104
rect 20477 -6165 20553 -6160
rect 21137 -2619 21213 -2614
rect 21137 -2675 21147 -2619
rect 21203 -2675 21213 -2619
rect 21137 -3819 21213 -2675
rect 21137 -3875 21147 -3819
rect 21203 -3875 21213 -3819
rect 21137 -5019 21213 -3875
rect 21137 -5075 21147 -5019
rect 21203 -5075 21213 -5019
rect 21137 -6219 21213 -5075
rect 21137 -6275 21147 -6219
rect 21203 -6275 21213 -6219
rect 21137 -6280 21213 -6275
rect 21336 -2766 21412 -2761
rect 21336 -2822 21346 -2766
rect 21402 -2822 21412 -2766
rect 21336 -3966 21412 -2822
rect 21336 -4022 21346 -3966
rect 21402 -4022 21412 -3966
rect 21336 -5166 21412 -4022
rect 21336 -5222 21346 -5166
rect 21402 -5222 21412 -5166
rect 21336 -6366 21412 -5222
rect 22256 -3204 22332 -2060
rect 22256 -3260 22266 -3204
rect 22322 -3260 22332 -3204
rect 22256 -4404 22332 -3260
rect 22256 -4460 22266 -4404
rect 22322 -4460 22332 -4404
rect 22256 -5604 22332 -4460
rect 22472 -3086 22548 -1942
rect 22472 -3142 22482 -3086
rect 22538 -3142 22548 -3086
rect 22472 -4286 22548 -3142
rect 22472 -4342 22482 -4286
rect 22538 -4342 22548 -4286
rect 22472 -5486 22548 -4342
rect 22472 -5542 22482 -5486
rect 22538 -5542 22548 -5486
rect 22472 -5547 22548 -5542
rect 22256 -5660 22266 -5604
rect 22322 -5660 22332 -5604
rect 22256 -5665 22332 -5660
rect 21336 -6422 21346 -6366
rect 21402 -6422 21412 -6366
rect 21336 -6427 21412 -6422
use sky130_fd_pr__nfet_g5v0d10v5_M9JYBS  sky130_fd_pr__nfet_g5v0d10v5_M9JYBS_0
array 0 4 1836 0 0 1000
timestamp 1711636687
transform 1 0 14305 0 1 -5938
box -118 -99 118 99
use sky130_fd_pr__nfet_g5v0d10v5_M9JYBS  sky130_fd_pr__nfet_g5v0d10v5_M9JYBS_1
array 0 4 1836 0 0 1000
timestamp 1711636687
transform -1 0 28993 0 1 -5938
box -118 -99 118 99
use sky130_fd_pr__nfet_g5v0d10v5_M9JYBS  sky130_fd_pr__nfet_g5v0d10v5_M9JYBS_2
array 0 4 1836 0 0 1000
timestamp 1711636687
transform 1 0 14305 0 1 -4738
box -118 -99 118 99
use sky130_fd_pr__nfet_g5v0d10v5_M9JYBS  sky130_fd_pr__nfet_g5v0d10v5_M9JYBS_3
array 0 4 1836 0 0 1000
timestamp 1711636687
transform -1 0 28993 0 1 -4738
box -118 -99 118 99
use sky130_fd_pr__nfet_g5v0d10v5_M9JYBS  sky130_fd_pr__nfet_g5v0d10v5_M9JYBS_4
array 0 4 1836 0 0 1000
timestamp 1711636687
transform 1 0 14305 0 1 -3538
box -118 -99 118 99
use sky130_fd_pr__nfet_g5v0d10v5_M9JYBS  sky130_fd_pr__nfet_g5v0d10v5_M9JYBS_5
array 0 4 1836 0 0 1000
timestamp 1711636687
transform -1 0 28993 0 1 -3538
box -118 -99 118 99
use sky130_fd_pr__nfet_g5v0d10v5_M9JYBS  sky130_fd_pr__nfet_g5v0d10v5_M9JYBS_6
array 0 4 1836 0 0 1000
timestamp 1711636687
transform 1 0 14305 0 1 -2338
box -118 -99 118 99
use sky130_fd_pr__nfet_g5v0d10v5_M9JYBS  sky130_fd_pr__nfet_g5v0d10v5_M9JYBS_7
array 0 4 1836 0 0 1000
timestamp 1711636687
transform -1 0 28993 0 1 -2338
box -118 -99 118 99
use sky130_fd_pr__nfet_g5v0d10v5_NXCGNM  sky130_fd_pr__nfet_g5v0d10v5_NXCGNM_0
array 0 4 1836 0 0 1000
timestamp 1711636687
transform 1 0 13387 0 1 -5938
box -858 -99 858 99
use sky130_fd_pr__nfet_g5v0d10v5_NXCGNM  sky130_fd_pr__nfet_g5v0d10v5_NXCGNM_1
array 0 4 1836 0 0 1000
timestamp 1711636687
transform 1 0 13387 0 1 -4738
box -858 -99 858 99
use sky130_fd_pr__nfet_g5v0d10v5_NXCGNM  sky130_fd_pr__nfet_g5v0d10v5_NXCGNM_2
array 0 4 1836 0 0 1000
timestamp 1711636687
transform -1 0 29911 0 1 -5938
box -858 -99 858 99
use sky130_fd_pr__nfet_g5v0d10v5_NXCGNM  sky130_fd_pr__nfet_g5v0d10v5_NXCGNM_3
array 0 4 1836 0 0 1000
timestamp 1711636687
transform -1 0 29911 0 1 -2338
box -858 -99 858 99
use sky130_fd_pr__nfet_g5v0d10v5_NXCGNM  sky130_fd_pr__nfet_g5v0d10v5_NXCGNM_4
array 0 4 1836 0 0 1000
timestamp 1711636687
transform 1 0 13387 0 1 -3538
box -858 -99 858 99
use sky130_fd_pr__nfet_g5v0d10v5_NXCGNM  sky130_fd_pr__nfet_g5v0d10v5_NXCGNM_5
array 0 4 1836 0 0 1000
timestamp 1711636687
transform -1 0 29911 0 1 -4738
box -858 -99 858 99
use sky130_fd_pr__nfet_g5v0d10v5_NXCGNM  sky130_fd_pr__nfet_g5v0d10v5_NXCGNM_6
array 0 4 1836 0 0 1000
timestamp 1711636687
transform 1 0 13387 0 1 -2338
box -858 -99 858 99
use sky130_fd_pr__nfet_g5v0d10v5_NXCGNM  sky130_fd_pr__nfet_g5v0d10v5_NXCGNM_7
array 0 4 1836 0 0 1000
timestamp 1711636687
transform -1 0 29911 0 1 -3538
box -858 -99 858 99
<< labels >>
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 ibias
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ena
port 3 nsew
rlabel metal3 22472 -5383 22472 -5383 1 vinp
port 5 n
rlabel metal3 22256 -5383 22256 -5383 1 vinn
port 4 n
rlabel metal1 11953 -1964 11953 -1964 1 avss
port 6 n
rlabel metal1 8329 -2444 8329 -2444 1 avdd
port 0 n
rlabel metal3 20477 -5367 20477 -5367 1 vt
port 7 n
rlabel metal3 21137 -5367 21137 -5367 1 vnn
rlabel metal3 21336 -5367 21336 -5367 1 vpp
<< end >>
