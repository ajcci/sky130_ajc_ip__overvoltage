magic
tech sky130A
magscale 1 2
timestamp 1712888861
<< error_p >>
rect 44483 16217 44557 16226
rect 44483 16161 44492 16217
rect 44483 16152 44557 16161
rect 44000 15969 44074 15978
rect 44483 15969 44557 15978
rect 44000 15913 44009 15969
rect 44483 15913 44492 15969
rect 44000 15904 44074 15913
rect 44483 15904 44557 15913
<< pwell >>
rect -2026 68336 42057 68472
rect -2026 38153 -1890 68336
rect 41921 38153 42057 68336
rect -2026 38017 42057 38153
<< psubdiff >>
rect -1990 68402 -1930 68436
rect 41961 68402 42021 68436
rect -1990 68376 -1956 68402
rect -1990 38087 -1956 38113
rect 41987 68376 42021 68402
rect 41987 38087 42021 38113
rect -1990 38053 -1930 38087
rect 41961 38053 42021 38087
<< psubdiffcont >>
rect -1930 68402 41961 68436
rect -1990 38113 -1956 68376
rect 41987 38113 42021 68376
rect -1930 38053 41961 38087
<< locali >>
rect -1990 68402 -1930 68436
rect 41961 68402 42021 68436
rect -1990 68376 -1956 68402
rect -1990 38087 -1956 38113
rect 41987 68376 42021 68402
rect 41987 38087 42021 38113
rect -1990 38053 -1930 38087
rect 41961 38053 42021 38087
rect 44279 16275 44407 16290
rect 44279 16177 44294 16275
rect 44392 16177 44407 16275
rect 44623 16275 44687 16290
rect 44279 16162 44407 16177
rect 44488 16206 44552 16221
rect 44488 16172 44503 16206
rect 44537 16172 44552 16206
rect 44488 16157 44552 16172
rect 44623 16177 44638 16275
rect 44672 16177 44687 16275
rect 44623 16162 44687 16177
rect 45359 16159 45417 16171
rect 45359 16125 45371 16159
rect 45405 16125 45417 16159
rect 45359 16113 45417 16125
rect 45203 16017 45331 16032
rect 45203 15919 45218 16017
rect 45316 15919 45331 16017
rect 45471 16017 45535 16032
rect 45203 15904 45331 15919
rect 45372 15953 45436 15968
rect 45372 15919 45387 15953
rect 45421 15919 45436 15953
rect 45372 15904 45436 15919
rect 45471 15919 45486 16017
rect 45520 15919 45535 16017
rect 45471 15904 45535 15919
rect 45317 15649 45445 15664
rect 45317 15615 45332 15649
rect 45430 15615 45445 15649
rect 45317 15600 45445 15615
<< viali >>
rect -1930 68402 41961 68436
rect -1990 38156 -1956 68349
rect 41987 38145 42021 68338
rect -1930 38053 41961 38087
rect 44294 16177 44392 16275
rect 44503 16172 44537 16206
rect 44638 16177 44672 16275
rect 45371 16125 45405 16159
rect 45218 15919 45316 16017
rect 45387 15919 45421 15953
rect 45486 15919 45520 16017
rect 45332 15615 45430 15649
rect 39436 15526 39484 15574
<< metal1 >>
rect -2030 68436 42061 68476
rect -2030 68402 -1930 68436
rect 41961 68402 42061 68436
rect -2030 68349 42061 68402
rect -2030 38156 -1990 68349
rect -1956 68338 42061 68349
rect -1956 68336 41987 68338
rect -1956 38156 -1890 68336
rect -2030 38153 -1890 38156
rect 41921 38153 41987 68336
rect -2030 38145 41987 38153
rect 42021 38145 42061 68338
rect -2030 38087 42061 38145
rect -2030 38053 -1930 38087
rect 41961 38053 42061 38087
rect -2030 38013 42061 38053
rect 573 27559 579 27959
rect 979 27559 985 27959
rect 44269 16289 44417 16300
rect 44269 16163 44280 16289
rect 44406 16163 44417 16289
rect 44618 16289 44692 16300
rect 44269 16152 44417 16163
rect 44483 16215 44557 16226
rect 44483 16163 44494 16215
rect 44546 16163 44557 16215
rect 44483 16152 44557 16163
rect 44618 16163 44629 16289
rect 44681 16163 44692 16289
rect 44618 16152 44692 16163
rect 45359 16159 45417 16171
rect 45359 16125 45371 16159
rect 45405 16125 45417 16159
rect 45359 16113 45417 16125
rect 44269 16041 44417 16052
rect 44269 15915 44280 16041
rect 44406 15915 44417 16041
rect 44618 16041 44692 16052
rect 44269 15904 44417 15915
rect 44483 15967 44557 15978
rect 44483 15915 44494 15967
rect 44546 15915 44557 15967
rect 44483 15904 44557 15915
rect 44618 15915 44629 16041
rect 44681 15915 44692 16041
rect 44618 15904 44692 15915
rect 44775 16026 44903 16032
rect 44775 15910 44781 16026
rect 44897 15910 44903 16026
rect 45043 16026 45107 16032
rect 44775 15904 44903 15910
rect 44944 15962 45008 15968
rect 44944 15910 44950 15962
rect 45002 15910 45008 15962
rect 44944 15904 45008 15910
rect 45043 15910 45049 16026
rect 45101 15910 45107 16026
rect 45043 15904 45107 15910
rect 45203 16026 45331 16032
rect 45203 15910 45209 16026
rect 45325 15910 45331 16026
rect 45471 16026 45535 16032
rect 45203 15904 45331 15910
rect 45372 15962 45436 15968
rect 45372 15910 45378 15962
rect 45430 15910 45436 15962
rect 45372 15904 45436 15910
rect 45471 15910 45477 16026
rect 45529 15910 45535 16026
rect 45471 15904 45535 15910
rect 38208 15800 38272 15806
rect 38208 15748 38214 15800
rect 38266 15748 38272 15800
rect 38208 15742 38272 15748
rect 38520 15799 38584 15805
rect 39151 15804 39215 15810
rect 38520 15747 38526 15799
rect 38578 15747 38584 15799
rect 38520 15741 38584 15747
rect 38835 15798 38899 15804
rect 38835 15746 38841 15798
rect 38893 15746 38899 15798
rect 39151 15752 39157 15804
rect 39209 15752 39215 15804
rect 39151 15746 39215 15752
rect 38835 15740 38899 15746
rect 45063 15732 45191 15738
rect 45063 15680 45069 15732
rect 45185 15680 45191 15732
rect 45063 15674 45191 15680
rect 45317 15658 45445 15664
rect 44627 15643 44775 15654
rect 38060 15580 38106 15612
rect 38376 15580 38422 15612
rect 38692 15580 38738 15612
rect 39008 15580 39054 15612
rect 39324 15580 39370 15612
rect 44627 15591 44638 15643
rect 44764 15591 44775 15643
rect 45317 15606 45323 15658
rect 45439 15606 45445 15658
rect 45317 15600 45445 15606
rect 39424 15580 39496 15587
rect 44627 15580 44775 15591
rect 38060 15534 38116 15580
rect 38208 15534 39430 15580
rect 39424 15520 39430 15534
rect 39490 15520 39496 15580
rect 39424 15513 39496 15520
rect 38495 11718 41643 12028
rect 41953 11718 41959 12028
rect 38553 11462 42086 11662
rect 42286 11462 42292 11662
rect 38481 11206 40724 11406
rect 40924 11206 40930 11406
<< via1 >>
rect 579 27559 979 27959
rect 44280 16275 44406 16289
rect 44280 16177 44294 16275
rect 44294 16177 44392 16275
rect 44392 16177 44406 16275
rect 44280 16163 44406 16177
rect 44494 16206 44546 16215
rect 44494 16172 44503 16206
rect 44503 16172 44537 16206
rect 44537 16172 44546 16206
rect 44494 16163 44546 16172
rect 44629 16275 44681 16289
rect 44629 16177 44638 16275
rect 44638 16177 44672 16275
rect 44672 16177 44681 16275
rect 44629 16163 44681 16177
rect 44280 15915 44406 16041
rect 44494 15915 44546 15967
rect 44629 15915 44681 16041
rect 44781 15910 44897 16026
rect 44950 15910 45002 15962
rect 45049 15910 45101 16026
rect 45209 16017 45325 16026
rect 45209 15919 45218 16017
rect 45218 15919 45316 16017
rect 45316 15919 45325 16017
rect 45209 15910 45325 15919
rect 45378 15953 45430 15962
rect 45378 15919 45387 15953
rect 45387 15919 45421 15953
rect 45421 15919 45430 15953
rect 45378 15910 45430 15919
rect 45477 16017 45529 16026
rect 45477 15919 45486 16017
rect 45486 15919 45520 16017
rect 45520 15919 45529 16017
rect 45477 15910 45529 15919
rect 38214 15748 38266 15800
rect 38526 15747 38578 15799
rect 38841 15746 38893 15798
rect 39157 15752 39209 15804
rect 45069 15680 45185 15732
rect 44638 15591 44764 15643
rect 45323 15649 45439 15658
rect 45323 15615 45332 15649
rect 45332 15615 45430 15649
rect 45430 15615 45439 15649
rect 45323 15606 45439 15615
rect 39430 15574 39490 15580
rect 39430 15526 39436 15574
rect 39436 15526 39484 15574
rect 39484 15526 39490 15574
rect 39430 15520 39490 15526
rect 41643 11718 41953 12028
rect 42086 11462 42286 11662
rect 40724 11206 40924 11406
<< metal2 >>
rect 579 27959 979 27965
rect 123 27494 523 27503
rect 123 25701 523 27094
rect 579 25705 979 27559
rect 8831 21182 8883 28879
rect 9797 21381 9857 28879
rect 10854 16753 10928 28879
rect 13054 13951 13118 28879
rect 25007 27689 25108 27698
rect 25007 26676 25108 27588
rect 40064 23473 40120 23480
rect 28660 23464 28724 23473
rect 22447 20766 22503 20773
rect 22445 20764 22505 20766
rect 22445 20708 22447 20764
rect 22503 20708 22505 20764
rect 20145 18358 20209 18362
rect 20140 18302 20149 18358
rect 20205 18302 20214 18358
rect 13054 13887 13154 13951
rect 13090 13778 13154 13887
rect 20145 13760 20209 18302
rect 20342 15399 20398 15406
rect 20340 15397 20400 15399
rect 20340 15341 20342 15397
rect 20398 15341 20400 15397
rect 20340 13974 20400 15341
rect 22445 13943 22505 20708
rect 24716 16553 24772 16560
rect 24714 16551 24774 16553
rect 24714 16495 24716 16551
rect 24772 16495 24774 16551
rect 24562 15905 24626 15914
rect 22612 15552 22668 15559
rect 22610 15550 22670 15552
rect 22610 15494 22612 15550
rect 22668 15494 22670 15550
rect 22610 13806 22670 15494
rect 24562 13881 24626 15841
rect 20145 13696 20396 13760
rect 20332 12238 20396 13696
rect 22453 13746 22670 13806
rect 24714 13765 24774 16495
rect 25935 16395 25991 18391
rect 26550 17837 26606 17842
rect 26546 17833 26610 17837
rect 26546 17777 26550 17833
rect 26606 17777 26610 17833
rect 25933 16386 25993 16395
rect 25933 16317 25993 16326
rect 26546 15049 26610 17777
rect 26693 17624 26749 17631
rect 26691 17622 26751 17624
rect 26691 17566 26693 17622
rect 26749 17566 26751 17622
rect 26691 15049 26751 17566
rect 28660 15726 28724 23400
rect 40062 23471 40122 23473
rect 40062 23415 40064 23471
rect 40120 23415 40122 23471
rect 39902 22793 39958 22800
rect 39900 22791 39960 22793
rect 28819 22772 28883 22781
rect 28819 15901 28883 22708
rect 39900 22735 39902 22791
rect 39958 22735 39960 22791
rect 39761 22113 39817 22120
rect 39759 22111 39819 22113
rect 29072 22093 29136 22102
rect 28941 21406 29005 21415
rect 28941 17842 29005 21342
rect 29072 18506 29136 22029
rect 39759 22055 39761 22111
rect 39817 22055 39819 22111
rect 39222 21433 39278 21440
rect 39220 21431 39280 21433
rect 39220 21375 39222 21431
rect 39278 21375 39280 21431
rect 32808 18510 32864 18515
rect 29072 18450 29076 18506
rect 29132 18450 29136 18506
rect 29072 18446 29136 18450
rect 32804 18506 32868 18510
rect 32804 18450 32808 18506
rect 32864 18450 32868 18506
rect 29076 18441 29132 18446
rect 28932 17837 29014 17842
rect 28932 17773 28941 17837
rect 29005 17773 29014 17837
rect 28932 17764 29014 17773
rect 31342 17765 31398 17772
rect 31340 17763 31400 17765
rect 31340 17707 31342 17763
rect 31398 17707 31400 17763
rect 28969 16005 29025 16012
rect 31340 16010 31400 17707
rect 31331 16005 31409 16010
rect 28819 15845 28823 15901
rect 28879 15845 28883 15901
rect 28819 15841 28883 15845
rect 28967 16003 29027 16005
rect 28967 15947 28969 16003
rect 29025 15947 29027 16003
rect 28823 15836 28879 15841
rect 28660 15670 28664 15726
rect 28720 15670 28724 15726
rect 28660 15666 28724 15670
rect 28664 15661 28720 15666
rect 28800 15263 28856 15270
rect 22453 12228 22513 13746
rect 24570 13705 24774 13765
rect 26541 14910 26610 15049
rect 26682 14952 26751 15049
rect 28798 15261 28858 15263
rect 28798 15205 28800 15261
rect 28856 15205 28858 15261
rect 28798 15049 28858 15205
rect 26541 13756 26605 14910
rect 26682 14012 26742 14952
rect 28798 14931 28859 15049
rect 28967 15044 29027 15947
rect 31331 15945 31340 16005
rect 31400 15945 31409 16005
rect 31331 15936 31409 15945
rect 30725 15730 30781 15735
rect 30915 15733 30971 15740
rect 30913 15731 30973 15733
rect 28799 13965 28859 14931
rect 28940 14928 29027 15044
rect 30721 15726 30785 15730
rect 30721 15670 30725 15726
rect 30781 15670 30785 15726
rect 30721 15049 30785 15670
rect 30913 15675 30915 15731
rect 30971 15675 30973 15731
rect 30913 15049 30973 15675
rect 32448 15561 32504 16631
rect 32446 15552 32506 15561
rect 32446 15483 32506 15492
rect 30721 14930 30786 15049
rect 28940 13780 29000 14928
rect 24570 12218 24630 13705
rect 26541 13692 26738 13756
rect 26674 12147 26738 13692
rect 28791 13720 29000 13780
rect 30722 13804 30786 14930
rect 30903 14925 30973 15049
rect 32804 15049 32868 18450
rect 33305 18200 33361 18207
rect 33303 18198 33363 18200
rect 33303 18142 33305 18198
rect 33361 18142 33363 18198
rect 33092 16562 33148 16631
rect 33090 16553 33150 16562
rect 33090 16484 33150 16493
rect 33303 15733 33363 18142
rect 34813 18069 34869 18076
rect 34811 18067 34871 18069
rect 34811 18011 34813 18067
rect 34869 18011 34871 18067
rect 33501 17904 33557 17911
rect 33303 15664 33363 15673
rect 33499 17902 33559 17904
rect 33499 17846 33501 17902
rect 33557 17846 33559 17902
rect 30903 13987 30963 14925
rect 32804 14887 32869 15049
rect 33013 15031 33073 15049
rect 32995 15022 33073 15031
rect 33051 14966 33073 15022
rect 32995 14957 33073 14966
rect 30722 13740 30962 13804
rect 28791 12233 28851 13720
rect 30898 12147 30962 13740
rect 32805 13753 32869 14887
rect 33013 13975 33073 14957
rect 33499 15024 33559 17846
rect 33736 15408 33792 16631
rect 33734 15399 33794 15408
rect 33734 15330 33794 15339
rect 34380 15272 34436 16631
rect 34378 15263 34438 15272
rect 34378 15194 34438 15203
rect 34811 15004 34871 18011
rect 39220 17909 39280 21375
rect 39363 20753 39419 20760
rect 39361 20751 39421 20753
rect 39361 20695 39363 20751
rect 39419 20695 39421 20751
rect 39361 18069 39421 20695
rect 39497 20071 39557 20073
rect 39490 20015 39499 20071
rect 39555 20015 39564 20071
rect 39497 19563 39557 20015
rect 39497 19503 39683 19563
rect 39497 19391 39561 19395
rect 39492 19335 39501 19391
rect 39557 19335 39566 19391
rect 39497 18362 39561 19335
rect 39497 18289 39561 18298
rect 39623 18200 39683 19503
rect 39623 18131 39683 18140
rect 39361 18000 39421 18009
rect 39211 17904 39289 17909
rect 39211 17844 39220 17904
rect 39280 17844 39289 17904
rect 39211 17835 39289 17844
rect 39759 17765 39819 22055
rect 39759 17696 39819 17705
rect 39900 17624 39960 22735
rect 39900 17555 39960 17564
rect 37727 17467 37783 17474
rect 40062 17467 40122 23415
rect 37725 17465 37785 17467
rect 37725 17409 37727 17465
rect 37783 17409 37785 17465
rect 36143 16877 36203 16886
rect 35024 15756 35080 16631
rect 35668 16004 35724 16640
rect 36143 16387 36203 16817
rect 36136 16331 36145 16387
rect 36201 16331 36210 16387
rect 36143 16329 36203 16331
rect 36312 16288 36368 16657
rect 36956 16570 37012 16647
rect 36954 16561 37014 16570
rect 36954 16492 37014 16501
rect 36310 16279 36370 16288
rect 36310 16210 36370 16219
rect 35666 15995 35726 16004
rect 35666 15926 35726 15935
rect 35022 15747 35082 15756
rect 35022 15678 35082 15687
rect 37725 15124 37785 17409
rect 40062 17398 40122 17407
rect 38201 16559 38275 16568
rect 38201 16503 38210 16559
rect 38266 16503 38275 16559
rect 38201 16498 38275 16503
rect 38208 15806 38268 16498
rect 44269 16291 44417 16300
rect 38528 16277 38588 16279
rect 38521 16221 38530 16277
rect 38586 16221 38595 16277
rect 38208 15800 38272 15806
rect 38528 15805 38588 16221
rect 44269 16161 44278 16291
rect 44408 16161 44417 16291
rect 44618 16291 44692 16300
rect 44269 16152 44417 16161
rect 44483 16217 44557 16226
rect 44483 16161 44492 16217
rect 44548 16161 44557 16217
rect 44483 16152 44557 16161
rect 44618 16161 44627 16291
rect 44683 16161 44692 16291
rect 44618 16152 44692 16161
rect 43785 16043 43933 16052
rect 38828 15993 38902 16002
rect 38828 15937 38837 15993
rect 38893 15937 38902 15993
rect 38828 15932 38902 15937
rect 38208 15748 38214 15800
rect 38266 15748 38272 15800
rect 38208 15742 38272 15748
rect 38520 15799 38588 15805
rect 38520 15747 38526 15799
rect 38578 15747 38588 15799
rect 38520 15745 38588 15747
rect 38835 15804 38895 15932
rect 43785 15913 43794 16043
rect 43924 15913 43933 16043
rect 44134 16043 44208 16052
rect 43785 15904 43933 15913
rect 44000 15969 44074 15978
rect 44000 15913 44009 15969
rect 44065 15913 44074 15969
rect 44000 15904 44074 15913
rect 44134 15913 44143 16043
rect 44199 15913 44208 16043
rect 44134 15904 44208 15913
rect 44269 16043 44417 16052
rect 44269 15913 44278 16043
rect 44408 15913 44417 16043
rect 44618 16043 44692 16052
rect 44269 15904 44417 15913
rect 44483 15969 44557 15978
rect 44483 15913 44492 15969
rect 44548 15913 44557 15969
rect 44483 15904 44557 15913
rect 44618 15913 44627 16043
rect 44683 15913 44692 16043
rect 44618 15904 44692 15913
rect 44775 16026 44903 16032
rect 44775 15910 44781 16026
rect 44897 15910 44903 16026
rect 45043 16026 45107 16032
rect 44775 15904 44903 15910
rect 44944 15962 45008 15968
rect 44944 15910 44950 15962
rect 45002 15910 45008 15962
rect 44944 15904 45008 15910
rect 45043 15910 45049 16026
rect 45101 15910 45107 16026
rect 45043 15904 45107 15910
rect 45203 16026 45331 16032
rect 45203 15910 45209 16026
rect 45325 15910 45331 16026
rect 45471 16026 45535 16032
rect 45203 15904 45331 15910
rect 45372 15962 45436 15968
rect 45372 15910 45378 15962
rect 45430 15910 45436 15962
rect 45372 15904 45436 15910
rect 45471 15910 45477 16026
rect 45529 15910 45535 16026
rect 45471 15904 45535 15910
rect 39149 15804 39216 15810
rect 38835 15798 38899 15804
rect 38835 15746 38841 15798
rect 38893 15746 38899 15798
rect 38520 15741 38584 15745
rect 38835 15740 38899 15746
rect 39149 15752 39157 15804
rect 39209 15752 39216 15804
rect 39149 15745 39216 15752
rect 39149 15689 39158 15745
rect 39214 15689 39223 15745
rect 45063 15732 45191 15738
rect 44143 15689 44291 15698
rect 39156 15687 39216 15689
rect 44143 15633 44152 15689
rect 44282 15633 44291 15689
rect 45063 15680 45069 15732
rect 45185 15680 45191 15732
rect 45063 15674 45191 15680
rect 45317 15658 45445 15664
rect 44143 15624 44291 15633
rect 44627 15645 44775 15654
rect 44627 15589 44636 15645
rect 44766 15589 44775 15645
rect 45317 15606 45323 15658
rect 45439 15606 45445 15658
rect 45317 15600 45445 15606
rect 39424 15580 39496 15587
rect 44627 15580 44775 15589
rect 39424 15520 39430 15580
rect 39490 15520 39496 15580
rect 39424 15513 39496 15520
rect 35330 15122 35390 15124
rect 35323 15066 35332 15122
rect 35388 15066 35397 15122
rect 35124 15011 35184 15049
rect 33499 14955 33559 14964
rect 34802 14944 34811 15004
rect 34871 14944 34880 15004
rect 35122 15002 35184 15011
rect 35178 14946 35184 15002
rect 35122 14937 35184 14946
rect 35124 13950 35184 14937
rect 35325 14932 35390 15066
rect 37725 15049 37785 15064
rect 35325 13812 35385 14932
rect 37225 13947 37307 13952
rect 37225 13883 37234 13947
rect 37298 13883 37307 13947
rect 37225 13875 37307 13883
rect 32805 13689 33074 13753
rect 33010 12151 33074 13689
rect 35131 13752 35385 13812
rect 35131 12271 35191 13752
rect 37225 12147 37234 12211
rect 37298 12147 37307 12211
rect 41632 12028 41964 12039
rect 41632 11718 41643 12028
rect 41953 11718 41964 12028
rect 41632 11707 41964 11718
rect 42077 11662 42295 11671
rect 42077 11462 42086 11662
rect 42286 11462 42295 11662
rect 42077 11453 42295 11462
rect 40715 11406 40933 11415
rect 40715 11206 40724 11406
rect 40924 11206 40933 11406
rect 40715 11197 40933 11206
rect 582 8086 972 8095
rect 582 7687 972 7696
rect 8809 -1091 9111 5783
rect 9164 -643 9466 5444
rect 9164 -954 9466 -945
rect 8809 -1402 9111 -1393
<< via2 >>
rect 123 27094 523 27494
rect 25007 27588 25108 27689
rect 28660 23400 28724 23464
rect 22447 20708 22503 20764
rect 20149 18302 20205 18358
rect 20342 15341 20398 15397
rect 24716 16495 24772 16551
rect 24562 15841 24626 15905
rect 22612 15494 22668 15550
rect 26550 17777 26606 17833
rect 25933 16326 25993 16386
rect 26693 17566 26749 17622
rect 40064 23415 40120 23471
rect 28819 22708 28883 22772
rect 39902 22735 39958 22791
rect 29072 22029 29136 22093
rect 28941 21342 29005 21406
rect 39761 22055 39817 22111
rect 39222 21375 39278 21431
rect 29076 18450 29132 18506
rect 32808 18450 32864 18506
rect 28941 17773 29005 17837
rect 31342 17707 31398 17763
rect 28823 15845 28879 15901
rect 28969 15947 29025 16003
rect 28664 15670 28720 15726
rect 28800 15205 28856 15261
rect 31340 15945 31400 16005
rect 30725 15670 30781 15726
rect 30915 15675 30971 15731
rect 32446 15492 32506 15552
rect 33305 18142 33361 18198
rect 33090 16493 33150 16553
rect 34813 18011 34869 18067
rect 33303 15673 33363 15733
rect 33501 17846 33557 17902
rect 32995 14966 33051 15022
rect 33734 15339 33794 15399
rect 34378 15203 34438 15263
rect 33499 14964 33559 15024
rect 39363 20695 39419 20751
rect 39499 20015 39555 20071
rect 39501 19335 39557 19391
rect 39497 18298 39561 18362
rect 39623 18140 39683 18200
rect 39361 18009 39421 18069
rect 39220 17844 39280 17904
rect 39759 17705 39819 17765
rect 39900 17564 39960 17624
rect 37727 17409 37783 17465
rect 36143 16817 36203 16877
rect 36145 16331 36201 16387
rect 36954 16501 37014 16561
rect 36310 16219 36370 16279
rect 35666 15935 35726 15995
rect 35022 15687 35082 15747
rect 40062 17407 40122 17467
rect 38210 16503 38266 16559
rect 38530 16221 38586 16277
rect 44278 16289 44408 16291
rect 44278 16163 44280 16289
rect 44280 16163 44406 16289
rect 44406 16163 44408 16289
rect 44278 16161 44408 16163
rect 44492 16215 44548 16217
rect 44492 16163 44494 16215
rect 44494 16163 44546 16215
rect 44546 16163 44548 16215
rect 44492 16161 44548 16163
rect 44627 16289 44683 16291
rect 44627 16163 44629 16289
rect 44629 16163 44681 16289
rect 44681 16163 44683 16289
rect 44627 16161 44683 16163
rect 38837 15937 38893 15993
rect 43794 15913 43924 16043
rect 44009 15913 44065 15969
rect 44143 15913 44199 16043
rect 44278 16041 44408 16043
rect 44278 15915 44280 16041
rect 44280 15915 44406 16041
rect 44406 15915 44408 16041
rect 44278 15913 44408 15915
rect 44492 15967 44548 15969
rect 44492 15915 44494 15967
rect 44494 15915 44546 15967
rect 44546 15915 44548 15967
rect 44492 15913 44548 15915
rect 44627 16041 44683 16043
rect 44627 15915 44629 16041
rect 44629 15915 44681 16041
rect 44681 15915 44683 16041
rect 44627 15913 44683 15915
rect 39158 15689 39214 15745
rect 44152 15633 44282 15689
rect 44636 15643 44766 15645
rect 44636 15591 44638 15643
rect 44638 15591 44764 15643
rect 44764 15591 44766 15643
rect 44636 15589 44766 15591
rect 39432 15522 39488 15578
rect 35332 15066 35388 15122
rect 34811 14944 34871 15004
rect 35122 14946 35178 15002
rect 37725 15064 37785 15124
rect 37234 13883 37298 13947
rect 37234 12147 37298 12211
rect 41643 11718 41953 12028
rect 42086 11462 42286 11662
rect 40724 11206 40924 11406
rect 582 7696 972 8086
rect 123 6835 523 7235
rect 9164 -945 9466 -643
rect 8809 -1393 9111 -1091
<< metal3 >>
rect -2433 28873 42464 28879
rect -2433 28485 -2427 28873
rect -2039 28806 42070 28873
rect -2039 28798 35511 28806
rect -2039 28485 30511 28798
rect -2433 28480 30511 28485
rect 30829 28488 35511 28798
rect 35829 28488 42070 28806
rect 30829 28485 42070 28488
rect 42458 28485 42464 28873
rect 30829 28480 42464 28485
rect -2433 28479 42464 28480
rect -2433 28413 42464 28419
rect -2433 28025 -1967 28413
rect -1579 28373 41610 28413
rect -1579 28055 31171 28373
rect 31489 28356 41610 28373
rect 31489 28055 36171 28356
rect -1579 28038 36171 28055
rect 36489 28038 41610 28356
rect -1579 28025 41610 28038
rect 41998 28025 42464 28413
rect -2433 28019 42464 28025
rect -2433 27953 42464 27959
rect -2433 27565 -1507 27953
rect -1119 27689 41150 27953
rect -1119 27588 25007 27689
rect 25108 27588 41150 27689
rect -1119 27565 41150 27588
rect 41538 27565 42464 27953
rect -2433 27559 42464 27565
rect -2433 27494 42464 27499
rect -2433 27493 123 27494
rect -2433 27105 -1047 27493
rect -659 27105 123 27493
rect -2433 27099 123 27105
rect 118 27094 123 27099
rect 523 27493 42464 27494
rect 523 27105 40690 27493
rect 41078 27105 42464 27493
rect 523 27099 42464 27105
rect 523 27094 528 27099
rect 118 27089 528 27094
rect 40059 23473 40125 23476
rect 39697 23471 40125 23473
rect 28655 23464 28729 23469
rect 28655 23400 28660 23464
rect 28724 23400 28729 23464
rect 39697 23415 40064 23471
rect 40120 23415 40125 23471
rect 39697 23413 40125 23415
rect 40059 23410 40125 23413
rect 28655 23395 28729 23400
rect 39897 22793 39963 22796
rect 39679 22791 39963 22793
rect 28814 22772 28888 22777
rect 28814 22708 28819 22772
rect 28883 22708 28888 22772
rect 39679 22735 39902 22791
rect 39958 22735 39963 22791
rect 39679 22733 39963 22735
rect 39897 22730 39963 22733
rect 28814 22703 28888 22708
rect 39756 22113 39822 22116
rect 39532 22111 39822 22113
rect 29067 22093 29141 22098
rect 29067 22029 29072 22093
rect 29136 22029 29141 22093
rect 39532 22055 39761 22111
rect 39817 22055 39822 22111
rect 39532 22053 39822 22055
rect 39756 22050 39822 22053
rect 29067 22024 29141 22029
rect 39217 21433 39283 21436
rect 39217 21431 39593 21433
rect 28936 21406 29010 21411
rect 28936 21342 28941 21406
rect 29005 21342 29010 21406
rect 39217 21375 39222 21431
rect 39278 21375 39593 21431
rect 39217 21373 39593 21375
rect 39217 21370 39283 21373
rect 28936 21337 29010 21342
rect 22442 20766 22508 20769
rect 22442 20764 28566 20766
rect 22442 20708 22447 20764
rect 22503 20708 28566 20764
rect 22442 20706 28566 20708
rect 39358 20753 39424 20756
rect 39358 20751 39731 20753
rect 22442 20703 22508 20706
rect 39358 20695 39363 20751
rect 39419 20695 39731 20751
rect 39358 20693 39731 20695
rect 39358 20690 39424 20693
rect 39494 20071 39560 20076
rect 39494 20015 39499 20071
rect 39555 20015 39560 20071
rect 39494 20010 39560 20015
rect 39496 19391 39562 19396
rect 39496 19335 39501 19391
rect 39557 19335 39562 19391
rect 39496 19330 39562 19335
rect 29071 18510 29137 18511
rect 32803 18510 32869 18511
rect 29071 18506 32869 18510
rect 29071 18450 29076 18506
rect 29132 18450 32808 18506
rect 32864 18450 32869 18506
rect 29071 18446 32869 18450
rect 29071 18445 29137 18446
rect 32803 18445 32869 18446
rect 20144 18362 20210 18363
rect 39492 18362 39566 18367
rect 20144 18358 39497 18362
rect 20144 18302 20149 18358
rect 20205 18302 39497 18358
rect 20144 18298 39497 18302
rect 39561 18298 39566 18362
rect 20144 18297 20210 18298
rect 39492 18293 39566 18298
rect 33300 18200 33366 18203
rect 39618 18200 39688 18205
rect 33300 18198 39623 18200
rect 33300 18142 33305 18198
rect 33361 18142 39623 18198
rect 33300 18140 39623 18142
rect 39683 18140 39688 18200
rect 33300 18137 33366 18140
rect 39618 18135 39688 18140
rect 34808 18069 34874 18072
rect 39356 18069 39426 18074
rect 34808 18067 39361 18069
rect 34808 18011 34813 18067
rect 34869 18011 39361 18067
rect 34808 18009 39361 18011
rect 39421 18009 39426 18069
rect 34808 18006 34874 18009
rect 39356 18004 39426 18009
rect 33496 17904 33562 17907
rect 39215 17904 39285 17909
rect 33496 17902 39220 17904
rect 33496 17846 33501 17902
rect 33557 17846 39220 17902
rect 33496 17844 39220 17846
rect 39280 17844 39285 17904
rect 26545 17837 26611 17838
rect 28936 17837 29010 17842
rect 33496 17841 33562 17844
rect 39215 17839 39285 17844
rect 26545 17833 28941 17837
rect 26545 17777 26550 17833
rect 26606 17777 28941 17833
rect 26545 17773 28941 17777
rect 29005 17773 29010 17837
rect 26545 17772 26611 17773
rect 28936 17768 29010 17773
rect 31337 17765 31403 17768
rect 39754 17765 39824 17770
rect 31337 17763 39759 17765
rect 31337 17707 31342 17763
rect 31398 17707 39759 17763
rect 31337 17705 39759 17707
rect 39819 17705 39824 17765
rect 31337 17702 31403 17705
rect 39754 17700 39824 17705
rect 26688 17624 26754 17627
rect 39895 17624 39965 17629
rect 26688 17622 39900 17624
rect 26688 17566 26693 17622
rect 26749 17566 39900 17622
rect 26688 17564 39900 17566
rect 39960 17564 39965 17624
rect 26688 17561 26754 17564
rect 39895 17559 39965 17564
rect 37722 17467 37788 17470
rect 40057 17467 40127 17472
rect 37722 17465 40062 17467
rect 37722 17409 37727 17465
rect 37783 17409 40062 17465
rect 37722 17407 40062 17409
rect 40122 17407 40127 17467
rect 37722 17404 37788 17407
rect 40057 17402 40127 17407
rect 36138 16877 36208 16882
rect 36138 16817 36143 16877
rect 36203 16817 42464 16877
rect 36138 16812 36208 16817
rect 36949 16561 37019 16566
rect 38205 16561 38271 16564
rect 24711 16553 24777 16556
rect 33085 16553 33155 16558
rect 24711 16551 33090 16553
rect 24711 16495 24716 16551
rect 24772 16495 33090 16551
rect 24711 16493 33090 16495
rect 33150 16493 33155 16553
rect 36949 16501 36954 16561
rect 37014 16559 42464 16561
rect 37014 16503 38210 16559
rect 38266 16503 42464 16559
rect 37014 16501 42464 16503
rect 36949 16496 37019 16501
rect 38205 16498 38271 16501
rect 24711 16490 24777 16493
rect 33085 16488 33155 16493
rect 25928 16386 25998 16391
rect 36140 16389 36206 16392
rect 28160 16387 36206 16389
rect 28160 16386 36145 16387
rect 25928 16326 25933 16386
rect 25993 16331 36145 16386
rect 36201 16331 36206 16387
rect 25993 16329 36206 16331
rect 25993 16326 28332 16329
rect 36140 16326 36206 16329
rect 25928 16321 25998 16326
rect 44269 16291 44417 16300
rect 36305 16279 36375 16284
rect 38525 16279 38591 16282
rect 36305 16219 36310 16279
rect 36370 16277 42464 16279
rect 36370 16221 38530 16277
rect 38586 16221 42464 16277
rect 36370 16219 42464 16221
rect 36305 16214 36375 16219
rect 38525 16216 38591 16219
rect 44269 16161 44278 16291
rect 44408 16161 44417 16291
rect 44618 16291 44692 16300
rect 44269 16152 44417 16161
rect 44483 16217 44557 16226
rect 44483 16161 44492 16217
rect 44548 16161 44557 16217
rect 44483 16152 44557 16161
rect 44618 16161 44627 16291
rect 44683 16161 44692 16291
rect 44618 16152 44692 16161
rect 43785 16043 43933 16052
rect 28964 16005 29030 16008
rect 31335 16005 31405 16010
rect 28964 16003 31340 16005
rect 28964 15947 28969 16003
rect 29025 15947 31340 16003
rect 28964 15945 31340 15947
rect 31400 15945 31405 16005
rect 28964 15942 29030 15945
rect 31335 15940 31405 15945
rect 35661 15995 35731 16000
rect 38832 15995 38898 15998
rect 35661 15935 35666 15995
rect 35726 15993 42464 15995
rect 35726 15937 38837 15993
rect 38893 15937 42464 15993
rect 35726 15935 42464 15937
rect 35661 15930 35731 15935
rect 38832 15932 38898 15935
rect 43785 15913 43794 16043
rect 43924 15913 43933 16043
rect 44134 16043 44208 16052
rect 24557 15905 24631 15910
rect 28818 15905 28884 15906
rect 24557 15841 24562 15905
rect 24626 15901 28884 15905
rect 43785 15904 43933 15913
rect 44000 15969 44074 15978
rect 44000 15913 44009 15969
rect 44065 15913 44074 15969
rect 44000 15904 44074 15913
rect 44134 15913 44143 16043
rect 44199 15913 44208 16043
rect 44134 15904 44208 15913
rect 44269 16043 44417 16052
rect 44269 15913 44278 16043
rect 44408 15913 44417 16043
rect 44618 16043 44692 16052
rect 44269 15904 44417 15913
rect 44483 15969 44557 15978
rect 44483 15913 44492 15969
rect 44548 15913 44557 15969
rect 44483 15904 44557 15913
rect 44618 15913 44627 16043
rect 44683 15913 44692 16043
rect 44618 15904 44692 15913
rect 24626 15845 28823 15901
rect 28879 15845 28884 15901
rect 24626 15841 28884 15845
rect 24557 15836 24631 15841
rect 28818 15840 28884 15841
rect 35017 15747 35087 15752
rect 39153 15747 39219 15750
rect 30910 15733 30976 15736
rect 33298 15733 33368 15738
rect 30910 15731 33303 15733
rect 28659 15730 28725 15731
rect 30720 15730 30786 15731
rect 28659 15726 30786 15730
rect 28659 15670 28664 15726
rect 28720 15670 30725 15726
rect 30781 15670 30786 15726
rect 30910 15675 30915 15731
rect 30971 15675 33303 15731
rect 30910 15673 33303 15675
rect 33363 15673 33368 15733
rect 35017 15687 35022 15747
rect 35082 15745 42464 15747
rect 35082 15689 39158 15745
rect 39214 15689 42464 15745
rect 35082 15687 42464 15689
rect 44143 15689 44291 15698
rect 35017 15682 35087 15687
rect 39153 15684 39219 15687
rect 30910 15670 30976 15673
rect 28659 15666 30786 15670
rect 33298 15668 33368 15673
rect 28659 15665 28725 15666
rect 30720 15665 30786 15666
rect 44143 15633 44152 15689
rect 44282 15633 44291 15689
rect 44143 15624 44291 15633
rect 44627 15645 44775 15654
rect 44627 15589 44636 15645
rect 44766 15589 44775 15645
rect 39427 15580 39493 15583
rect 41626 15580 41632 15582
rect 39427 15578 41632 15580
rect 22607 15552 22673 15555
rect 32441 15552 32511 15557
rect 22607 15550 32446 15552
rect 22607 15494 22612 15550
rect 22668 15494 32446 15550
rect 22607 15492 32446 15494
rect 32506 15492 32511 15552
rect 39427 15522 39432 15578
rect 39488 15522 41632 15578
rect 39427 15520 41632 15522
rect 39427 15517 39493 15520
rect 41626 15518 41632 15520
rect 41696 15518 41702 15582
rect 44627 15580 44775 15589
rect 22607 15489 22673 15492
rect 32441 15487 32511 15492
rect 20337 15399 20403 15402
rect 33729 15399 33799 15404
rect 20337 15397 33734 15399
rect 20337 15341 20342 15397
rect 20398 15341 33734 15397
rect 20337 15339 33734 15341
rect 33794 15339 33799 15399
rect 20337 15336 20403 15339
rect 33729 15334 33799 15339
rect 28795 15263 28861 15266
rect 34373 15263 34443 15268
rect 28795 15261 34378 15263
rect 28795 15205 28800 15261
rect 28856 15205 34378 15261
rect 28795 15203 34378 15205
rect 34438 15203 34443 15263
rect 28795 15200 28861 15203
rect 34373 15198 34443 15203
rect 35327 15124 35393 15127
rect 37720 15124 37790 15129
rect 35327 15122 37725 15124
rect 35327 15066 35332 15122
rect 35388 15066 37725 15122
rect 35327 15064 37725 15066
rect 37785 15064 37790 15124
rect 35327 15061 35393 15064
rect 37720 15059 37790 15064
rect 32990 15024 33056 15027
rect 33494 15024 33564 15029
rect 32990 15022 33499 15024
rect 32990 14966 32995 15022
rect 33051 14966 33499 15022
rect 32990 14964 33499 14966
rect 33559 14964 33564 15024
rect 32990 14961 33056 14964
rect 33494 14959 33564 14964
rect 34806 15004 34876 15009
rect 35117 15004 35183 15007
rect 34806 14944 34811 15004
rect 34871 15002 35183 15004
rect 34871 14946 35122 15002
rect 35178 14946 35183 15002
rect 34871 14944 35183 14946
rect 34806 14939 34876 14944
rect 35117 14941 35183 14944
rect 4513 14168 4583 14238
rect 37229 13947 37303 13952
rect 37229 13883 37234 13947
rect 37298 13883 42464 13947
rect 37229 13878 37303 13883
rect 37229 12211 37303 12216
rect 37229 12147 37234 12211
rect 37298 12147 42464 12211
rect 37229 12142 37303 12147
rect 41632 12033 41964 12039
rect 41632 11713 41638 12033
rect 41958 11713 41964 12033
rect 41632 11707 41964 11713
rect 42077 11662 42295 11671
rect 42077 11462 42086 11662
rect 42286 11462 42295 11662
rect 42077 11453 42295 11462
rect 40715 11406 40933 11415
rect 40715 11206 40724 11406
rect 40924 11206 40933 11406
rect 40715 11197 40933 11206
rect -1518 8091 -1113 8096
rect -1518 8090 977 8091
rect -1518 7692 -1512 8090
rect -1114 8086 977 8090
rect -1114 7696 582 8086
rect 972 7696 977 8086
rect -1114 7692 977 7696
rect -1518 7691 977 7692
rect -1518 7686 -1113 7691
rect 118 7235 528 7240
rect -1056 6835 -1050 7235
rect -650 6835 123 7235
rect 523 6835 528 7235
rect 118 6830 528 6835
rect -2433 -616 42464 -610
rect -2433 -1004 -1047 -616
rect -659 -643 40690 -616
rect -659 -945 9164 -643
rect 9466 -945 40690 -643
rect -659 -1004 40690 -945
rect 41078 -1004 42464 -616
rect -2433 -1010 42464 -1004
rect -2433 -1076 42464 -1070
rect -2433 -1464 -1507 -1076
rect -1119 -1091 41150 -1076
rect -1119 -1393 8809 -1091
rect 9111 -1393 41150 -1091
rect -1119 -1464 41150 -1393
rect 41538 -1464 42464 -1076
rect -2433 -1470 42464 -1464
rect -2433 -1536 42464 -1530
rect -2433 -1924 -1967 -1536
rect -1579 -1924 41610 -1536
rect 41998 -1924 42464 -1536
rect -2433 -1930 42464 -1924
rect -2433 -1996 42464 -1990
rect -2433 -2384 -2427 -1996
rect -2039 -2384 42070 -1996
rect 42458 -2384 42464 -1996
rect -2433 -2390 42464 -2384
<< via3 >>
rect -2427 28485 -2039 28873
rect 30511 28480 30829 28798
rect 35511 28488 35829 28806
rect 42070 28485 42458 28873
rect -1967 28025 -1579 28413
rect 31171 28055 31489 28373
rect 36171 28038 36489 28356
rect 41610 28025 41998 28413
rect -1507 27565 -1119 27953
rect 41150 27565 41538 27953
rect -1047 27105 -659 27493
rect 40690 27105 41078 27493
rect 41632 15518 41696 15582
rect 41638 12028 41958 12033
rect 41638 11718 41643 12028
rect 41643 11718 41953 12028
rect 41953 11718 41958 12028
rect 41638 11713 41958 11718
rect 42086 11462 42286 11662
rect 40724 11206 40924 11406
rect -1512 7692 -1114 8090
rect -1050 6835 -650 7235
rect -1047 -1004 -659 -616
rect 40690 -1004 41078 -616
rect -1507 -1464 -1119 -1076
rect 41150 -1464 41538 -1076
rect -1967 -1924 -1579 -1536
rect 41610 -1924 41998 -1536
rect -2427 -2384 -2039 -1996
rect 42070 -2384 42458 -1996
<< metal4 >>
rect -2433 28873 -2033 28880
rect -2433 28485 -2427 28873
rect -2039 28485 -2033 28873
rect -2433 -1996 -2033 28485
rect -2433 -2384 -2427 -1996
rect -2039 -2384 -2033 -1996
rect -2433 -2390 -2033 -2384
rect -1973 28413 -1573 28880
rect -1973 28025 -1967 28413
rect -1579 28025 -1573 28413
rect -1973 -1536 -1573 28025
rect -1973 -1924 -1967 -1536
rect -1579 -1924 -1573 -1536
rect -1973 -2390 -1573 -1924
rect -1513 27953 -1113 28880
rect -1513 27565 -1507 27953
rect -1119 27565 -1113 27953
rect -1513 8090 -1113 27565
rect -1513 7692 -1512 8090
rect -1114 7692 -1113 8090
rect -1513 -1076 -1113 7692
rect -1513 -1464 -1507 -1076
rect -1119 -1464 -1113 -1076
rect -1513 -2390 -1113 -1464
rect -1053 27493 -653 28880
rect 35510 28806 35830 28807
rect -1053 27105 -1047 27493
rect -659 27105 -653 27493
rect -1053 7236 -653 27105
rect 30510 28798 30830 28799
rect 30510 28480 30511 28798
rect 30829 28480 30830 28798
rect 30510 26029 30830 28480
rect 35510 28488 35511 28806
rect 35829 28488 35830 28806
rect 31170 28373 31490 28374
rect 31170 28055 31171 28373
rect 31489 28055 31490 28373
rect 31170 25980 31490 28055
rect 35510 26095 35830 28488
rect 36170 28356 36490 28357
rect 36170 28038 36171 28356
rect 36489 28038 36490 28356
rect 36170 26015 36490 28038
rect 40684 27493 41084 28880
rect 40684 27105 40690 27493
rect 41078 27105 41084 27493
rect 40684 11406 41084 27105
rect 40684 11206 40724 11406
rect 40924 11206 41084 11406
rect -1053 7235 -649 7236
rect -1053 6835 -1050 7235
rect -650 6835 -649 7235
rect -1053 6834 -649 6835
rect -1053 -616 -653 6834
rect -1053 -1004 -1047 -616
rect -659 -1004 -653 -616
rect -1053 -2390 -653 -1004
rect 40684 -616 41084 11206
rect 40684 -1004 40690 -616
rect 41078 -1004 41084 -616
rect 40684 -2390 41084 -1004
rect 41144 27953 41544 28880
rect 41144 27565 41150 27953
rect 41538 27565 41544 27953
rect 41144 -1076 41544 27565
rect 41144 -1464 41150 -1076
rect 41538 -1464 41544 -1076
rect 41144 -2390 41544 -1464
rect 41604 28413 42004 28880
rect 41604 28025 41610 28413
rect 41998 28025 42004 28413
rect 41604 20547 42004 28025
rect 41604 20275 41689 20547
rect 41961 20275 42004 20547
rect 41604 15582 42004 20275
rect 41604 15518 41632 15582
rect 41696 15518 42004 15582
rect 41604 12033 42004 15518
rect 41604 11713 41638 12033
rect 41958 11713 42004 12033
rect 41604 -1536 42004 11713
rect 41604 -1924 41610 -1536
rect 41998 -1924 42004 -1536
rect 41604 -2390 42004 -1924
rect 42064 28873 42464 28880
rect 42064 28485 42070 28873
rect 42458 28485 42464 28873
rect 42064 19887 42464 28485
rect 42064 19615 42146 19887
rect 42418 19615 42464 19887
rect 42064 11662 42464 19615
rect 42064 11462 42086 11662
rect 42286 11462 42464 11662
rect 42064 -1996 42464 11462
rect 42064 -2384 42070 -1996
rect 42458 -2384 42464 -1996
rect 42064 -2390 42464 -2384
<< via4 >>
rect 41689 20275 41961 20547
rect 42146 19615 42418 19887
<< metal5 >>
rect 38371 20547 41985 20571
rect 38371 20275 41689 20547
rect 41961 20275 41985 20547
rect 38371 20251 41985 20275
rect 38371 19887 42442 19911
rect 38371 19615 42146 19887
rect 42418 19615 42442 19887
rect 38371 19591 42442 19615
use overvoltage_ana  overvoltage_ana_0
timestamp 1712718737
transform 1 0 28385 0 1 16000
box -29038 -16610 12299 11100
use overvoltage_dig  overvoltage_dig_0
timestamp 1712531369
transform 1 0 28566 0 1 16575
box 0 0 12000 9840
use sky130_fd_pr__nfet_01v8_9UEC9F  sky130_fd_pr__nfet_01v8_9UEC9F_0
timestamp 1712887115
transform 1 0 38715 0 1 15712
box -799 -310 799 310
<< labels >>
flabel metal3 894 -1930 894 -1930 0 FreeSans 1600 0 0 0 dvss
port 4 nsew
flabel metal3 894 -1470 894 -1470 0 FreeSans 1600 0 0 0 avss
port 2 nsew
flabel metal3 894 -1010 894 -1010 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal3 42464 15715 42464 15715 0 FreeSans 1280 0 0 0 otrip[0]
port 11 nsew
flabel metal3 42464 15964 42464 15964 0 FreeSans 1280 0 0 0 otrip[1]
port 10 nsew
flabel metal3 42464 16248 42464 16248 0 FreeSans 1280 0 0 0 otrip[2]
port 9 nsew
flabel metal3 42464 16529 42464 16529 0 FreeSans 1280 0 0 0 otrip[3]
port 8 nsew
flabel metal3 42464 16846 42464 16846 0 FreeSans 1280 0 0 0 ovout
port 6 nsew
flabel metal2 10891 28879 10891 28879 0 FreeSans 1280 0 0 0 itest
port 7 nsew
flabel metal2 8857 28879 8857 28879 0 FreeSans 1280 0 0 0 vbg_1v2
port 5 nsew
flabel metal2 9828 28879 9828 28879 0 FreeSans 1280 0 0 0 vin
port 12 nsew
flabel metal3 42464 12177 42464 12177 0 FreeSans 1280 0 0 0 ena
port 13 nsew
flabel metal3 42464 13915 42464 13915 0 FreeSans 1280 0 0 0 isrc_sel
port 14 nsew
flabel metal2 13085 28879 13085 28879 0 FreeSans 1280 0 0 0 ibg_200n
port 15 nsew
flabel metal3 894 -2390 894 -2390 0 FreeSans 1600 0 0 0 dvdd
port 3 nsew
<< end >>
