*This is the extracted netlist from layout

.subckt sky130_ajc_ip__overvoltage dvdd dvss otrip otrip_decoded

*Digital route extracted from layout
xIdig dvdd dvss otrip otrip_decoded overvoltage_dig

.ends

.subckt overvoltage_dig VPWR VGND otrip otrip_decoded
xbuf2 otrip VGND VGND VPWR VPWR otrip_decoded sky130_fd_sc_hd__buf_2
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
