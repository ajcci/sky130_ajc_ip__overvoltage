magic
tech sky130A
magscale 1 2
timestamp 1712027638
<< nwell >>
rect -1841 -4145 1841 4145
<< mvnsubdiff >>
rect -1775 4067 1775 4079
rect -1775 4033 -1667 4067
rect 1667 4033 1775 4067
rect -1775 4021 1775 4033
rect -1775 3971 -1717 4021
rect -1775 -3971 -1763 3971
rect -1729 -3971 -1717 3971
rect 1717 3971 1775 4021
rect -1775 -4021 -1717 -3971
rect 1717 -3971 1729 3971
rect 1763 -3971 1775 3971
rect 1717 -4021 1775 -3971
rect -1775 -4033 1775 -4021
rect -1775 -4067 -1667 -4033
rect 1667 -4067 1775 -4033
rect -1775 -4079 1775 -4067
<< mvnsubdiffcont >>
rect -1667 4033 1667 4067
rect -1763 -3971 -1729 3971
rect 1729 -3971 1763 3971
rect -1667 -4067 1667 -4033
<< xpolycontact >>
rect -1612 3484 -1542 3916
rect -1612 -3916 -1542 -3484
rect -1446 3484 -1376 3916
rect -1446 -3916 -1376 -3484
rect -1280 3484 -1210 3916
rect -1280 -3916 -1210 -3484
rect -1114 3484 -1044 3916
rect -1114 -3916 -1044 -3484
rect -948 3484 -878 3916
rect -948 -3916 -878 -3484
rect -782 3484 -712 3916
rect -782 -3916 -712 -3484
rect -616 3484 -546 3916
rect -616 -3916 -546 -3484
rect -450 3484 -380 3916
rect -450 -3916 -380 -3484
rect -284 3484 -214 3916
rect -284 -3916 -214 -3484
rect -118 3484 -48 3916
rect -118 -3916 -48 -3484
rect 48 3484 118 3916
rect 48 -3916 118 -3484
rect 214 3484 284 3916
rect 214 -3916 284 -3484
rect 380 3484 450 3916
rect 380 -3916 450 -3484
rect 546 3484 616 3916
rect 546 -3916 616 -3484
rect 712 3484 782 3916
rect 712 -3916 782 -3484
rect 878 3484 948 3916
rect 878 -3916 948 -3484
rect 1044 3484 1114 3916
rect 1044 -3916 1114 -3484
rect 1210 3484 1280 3916
rect 1210 -3916 1280 -3484
rect 1376 3484 1446 3916
rect 1376 -3916 1446 -3484
rect 1542 3484 1612 3916
rect 1542 -3916 1612 -3484
<< xpolyres >>
rect -1612 -3484 -1542 3484
rect -1446 -3484 -1376 3484
rect -1280 -3484 -1210 3484
rect -1114 -3484 -1044 3484
rect -948 -3484 -878 3484
rect -782 -3484 -712 3484
rect -616 -3484 -546 3484
rect -450 -3484 -380 3484
rect -284 -3484 -214 3484
rect -118 -3484 -48 3484
rect 48 -3484 118 3484
rect 214 -3484 284 3484
rect 380 -3484 450 3484
rect 546 -3484 616 3484
rect 712 -3484 782 3484
rect 878 -3484 948 3484
rect 1044 -3484 1114 3484
rect 1210 -3484 1280 3484
rect 1376 -3484 1446 3484
rect 1542 -3484 1612 3484
<< locali >>
rect -1763 4033 -1667 4067
rect 1667 4033 1763 4067
rect -1763 3971 -1729 4033
rect 1729 3971 1763 4033
rect -1763 -4033 -1729 -3971
rect 1729 -4033 1763 -3971
rect -1763 -4067 -1667 -4033
rect 1667 -4067 1763 -4033
<< viali >>
rect -1596 3501 -1558 3898
rect -1430 3501 -1392 3898
rect -1264 3501 -1226 3898
rect -1098 3501 -1060 3898
rect -932 3501 -894 3898
rect -766 3501 -728 3898
rect -600 3501 -562 3898
rect -434 3501 -396 3898
rect -268 3501 -230 3898
rect -102 3501 -64 3898
rect 64 3501 102 3898
rect 230 3501 268 3898
rect 396 3501 434 3898
rect 562 3501 600 3898
rect 728 3501 766 3898
rect 894 3501 932 3898
rect 1060 3501 1098 3898
rect 1226 3501 1264 3898
rect 1392 3501 1430 3898
rect 1558 3501 1596 3898
rect -1596 -3898 -1558 -3501
rect -1430 -3898 -1392 -3501
rect -1264 -3898 -1226 -3501
rect -1098 -3898 -1060 -3501
rect -932 -3898 -894 -3501
rect -766 -3898 -728 -3501
rect -600 -3898 -562 -3501
rect -434 -3898 -396 -3501
rect -268 -3898 -230 -3501
rect -102 -3898 -64 -3501
rect 64 -3898 102 -3501
rect 230 -3898 268 -3501
rect 396 -3898 434 -3501
rect 562 -3898 600 -3501
rect 728 -3898 766 -3501
rect 894 -3898 932 -3501
rect 1060 -3898 1098 -3501
rect 1226 -3898 1264 -3501
rect 1392 -3898 1430 -3501
rect 1558 -3898 1596 -3501
<< metal1 >>
rect -1602 3898 -1552 3910
rect -1602 3501 -1596 3898
rect -1558 3501 -1552 3898
rect -1602 3489 -1552 3501
rect -1436 3898 -1386 3910
rect -1436 3501 -1430 3898
rect -1392 3501 -1386 3898
rect -1436 3489 -1386 3501
rect -1270 3898 -1220 3910
rect -1270 3501 -1264 3898
rect -1226 3501 -1220 3898
rect -1270 3489 -1220 3501
rect -1104 3898 -1054 3910
rect -1104 3501 -1098 3898
rect -1060 3501 -1054 3898
rect -1104 3489 -1054 3501
rect -938 3898 -888 3910
rect -938 3501 -932 3898
rect -894 3501 -888 3898
rect -938 3489 -888 3501
rect -772 3898 -722 3910
rect -772 3501 -766 3898
rect -728 3501 -722 3898
rect -772 3489 -722 3501
rect -606 3898 -556 3910
rect -606 3501 -600 3898
rect -562 3501 -556 3898
rect -606 3489 -556 3501
rect -440 3898 -390 3910
rect -440 3501 -434 3898
rect -396 3501 -390 3898
rect -440 3489 -390 3501
rect -274 3898 -224 3910
rect -274 3501 -268 3898
rect -230 3501 -224 3898
rect -274 3489 -224 3501
rect -108 3898 -58 3910
rect -108 3501 -102 3898
rect -64 3501 -58 3898
rect -108 3489 -58 3501
rect 58 3898 108 3910
rect 58 3501 64 3898
rect 102 3501 108 3898
rect 58 3489 108 3501
rect 224 3898 274 3910
rect 224 3501 230 3898
rect 268 3501 274 3898
rect 224 3489 274 3501
rect 390 3898 440 3910
rect 390 3501 396 3898
rect 434 3501 440 3898
rect 390 3489 440 3501
rect 556 3898 606 3910
rect 556 3501 562 3898
rect 600 3501 606 3898
rect 556 3489 606 3501
rect 722 3898 772 3910
rect 722 3501 728 3898
rect 766 3501 772 3898
rect 722 3489 772 3501
rect 888 3898 938 3910
rect 888 3501 894 3898
rect 932 3501 938 3898
rect 888 3489 938 3501
rect 1054 3898 1104 3910
rect 1054 3501 1060 3898
rect 1098 3501 1104 3898
rect 1054 3489 1104 3501
rect 1220 3898 1270 3910
rect 1220 3501 1226 3898
rect 1264 3501 1270 3898
rect 1220 3489 1270 3501
rect 1386 3898 1436 3910
rect 1386 3501 1392 3898
rect 1430 3501 1436 3898
rect 1386 3489 1436 3501
rect 1552 3898 1602 3910
rect 1552 3501 1558 3898
rect 1596 3501 1602 3898
rect 1552 3489 1602 3501
rect -1602 -3501 -1552 -3489
rect -1602 -3898 -1596 -3501
rect -1558 -3898 -1552 -3501
rect -1602 -3910 -1552 -3898
rect -1436 -3501 -1386 -3489
rect -1436 -3898 -1430 -3501
rect -1392 -3898 -1386 -3501
rect -1436 -3910 -1386 -3898
rect -1270 -3501 -1220 -3489
rect -1270 -3898 -1264 -3501
rect -1226 -3898 -1220 -3501
rect -1270 -3910 -1220 -3898
rect -1104 -3501 -1054 -3489
rect -1104 -3898 -1098 -3501
rect -1060 -3898 -1054 -3501
rect -1104 -3910 -1054 -3898
rect -938 -3501 -888 -3489
rect -938 -3898 -932 -3501
rect -894 -3898 -888 -3501
rect -938 -3910 -888 -3898
rect -772 -3501 -722 -3489
rect -772 -3898 -766 -3501
rect -728 -3898 -722 -3501
rect -772 -3910 -722 -3898
rect -606 -3501 -556 -3489
rect -606 -3898 -600 -3501
rect -562 -3898 -556 -3501
rect -606 -3910 -556 -3898
rect -440 -3501 -390 -3489
rect -440 -3898 -434 -3501
rect -396 -3898 -390 -3501
rect -440 -3910 -390 -3898
rect -274 -3501 -224 -3489
rect -274 -3898 -268 -3501
rect -230 -3898 -224 -3501
rect -274 -3910 -224 -3898
rect -108 -3501 -58 -3489
rect -108 -3898 -102 -3501
rect -64 -3898 -58 -3501
rect -108 -3910 -58 -3898
rect 58 -3501 108 -3489
rect 58 -3898 64 -3501
rect 102 -3898 108 -3501
rect 58 -3910 108 -3898
rect 224 -3501 274 -3489
rect 224 -3898 230 -3501
rect 268 -3898 274 -3501
rect 224 -3910 274 -3898
rect 390 -3501 440 -3489
rect 390 -3898 396 -3501
rect 434 -3898 440 -3501
rect 390 -3910 440 -3898
rect 556 -3501 606 -3489
rect 556 -3898 562 -3501
rect 600 -3898 606 -3501
rect 556 -3910 606 -3898
rect 722 -3501 772 -3489
rect 722 -3898 728 -3501
rect 766 -3898 772 -3501
rect 722 -3910 772 -3898
rect 888 -3501 938 -3489
rect 888 -3898 894 -3501
rect 932 -3898 938 -3501
rect 888 -3910 938 -3898
rect 1054 -3501 1104 -3489
rect 1054 -3898 1060 -3501
rect 1098 -3898 1104 -3501
rect 1054 -3910 1104 -3898
rect 1220 -3501 1270 -3489
rect 1220 -3898 1226 -3501
rect 1264 -3898 1270 -3501
rect 1220 -3910 1270 -3898
rect 1386 -3501 1436 -3489
rect 1386 -3898 1392 -3501
rect 1430 -3898 1436 -3501
rect 1386 -3910 1436 -3898
rect 1552 -3501 1602 -3489
rect 1552 -3898 1558 -3501
rect 1596 -3898 1602 -3501
rect 1552 -3910 1602 -3898
<< properties >>
string FIXED_BBOX -1746 -4050 1746 4050
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 0.350 l 35 m 1 nx 20 wmin 0.350 lmin 0.50 rho 2000 val 201.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 1 hv_guard 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
