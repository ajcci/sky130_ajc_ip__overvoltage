magic
tech sky130A
timestamp 1712109191
<< pwell >>
rect -1601 -379 1601 379
<< mvnmos >>
rect -1487 -250 -1087 250
rect -1058 -250 -658 250
rect -629 -250 -229 250
rect -200 -250 200 250
rect 229 -250 629 250
rect 658 -250 1058 250
rect 1087 -250 1487 250
<< mvndiff >>
rect -1516 244 -1487 250
rect -1516 -244 -1510 244
rect -1493 -244 -1487 244
rect -1516 -250 -1487 -244
rect -1087 244 -1058 250
rect -1087 -244 -1081 244
rect -1064 -244 -1058 244
rect -1087 -250 -1058 -244
rect -658 244 -629 250
rect -658 -244 -652 244
rect -635 -244 -629 244
rect -658 -250 -629 -244
rect -229 244 -200 250
rect -229 -244 -223 244
rect -206 -244 -200 244
rect -229 -250 -200 -244
rect 200 244 229 250
rect 200 -244 206 244
rect 223 -244 229 244
rect 200 -250 229 -244
rect 629 244 658 250
rect 629 -244 635 244
rect 652 -244 658 244
rect 629 -250 658 -244
rect 1058 244 1087 250
rect 1058 -244 1064 244
rect 1081 -244 1087 244
rect 1058 -250 1087 -244
rect 1487 244 1516 250
rect 1487 -244 1493 244
rect 1510 -244 1516 244
rect 1487 -250 1516 -244
<< mvndiffc >>
rect -1510 -244 -1493 244
rect -1081 -244 -1064 244
rect -652 -244 -635 244
rect -223 -244 -206 244
rect 206 -244 223 244
rect 635 -244 652 244
rect 1064 -244 1081 244
rect 1493 -244 1510 244
<< mvpsubdiff >>
rect -1583 355 1583 361
rect -1583 338 -1529 355
rect 1529 338 1583 355
rect -1583 332 1583 338
rect -1583 307 -1554 332
rect -1583 -307 -1577 307
rect -1560 -307 -1554 307
rect 1554 307 1583 332
rect -1583 -332 -1554 -307
rect 1554 -307 1560 307
rect 1577 -307 1583 307
rect 1554 -332 1583 -307
rect -1583 -338 1583 -332
rect -1583 -355 -1529 -338
rect 1529 -355 1583 -338
rect -1583 -361 1583 -355
<< mvpsubdiffcont >>
rect -1529 338 1529 355
rect -1577 -307 -1560 307
rect 1560 -307 1577 307
rect -1529 -355 1529 -338
<< poly >>
rect -1487 286 -1087 294
rect -1487 269 -1479 286
rect -1095 269 -1087 286
rect -1487 250 -1087 269
rect -1058 286 -658 294
rect -1058 269 -1050 286
rect -666 269 -658 286
rect -1058 250 -658 269
rect -629 286 -229 294
rect -629 269 -621 286
rect -237 269 -229 286
rect -629 250 -229 269
rect -200 286 200 294
rect -200 269 -192 286
rect 192 269 200 286
rect -200 250 200 269
rect 229 286 629 294
rect 229 269 237 286
rect 621 269 629 286
rect 229 250 629 269
rect 658 286 1058 294
rect 658 269 666 286
rect 1050 269 1058 286
rect 658 250 1058 269
rect 1087 286 1487 294
rect 1087 269 1095 286
rect 1479 269 1487 286
rect 1087 250 1487 269
rect -1487 -269 -1087 -250
rect -1487 -286 -1479 -269
rect -1095 -286 -1087 -269
rect -1487 -294 -1087 -286
rect -1058 -269 -658 -250
rect -1058 -286 -1050 -269
rect -666 -286 -658 -269
rect -1058 -294 -658 -286
rect -629 -269 -229 -250
rect -629 -286 -621 -269
rect -237 -286 -229 -269
rect -629 -294 -229 -286
rect -200 -269 200 -250
rect -200 -286 -192 -269
rect 192 -286 200 -269
rect -200 -294 200 -286
rect 229 -269 629 -250
rect 229 -286 237 -269
rect 621 -286 629 -269
rect 229 -294 629 -286
rect 658 -269 1058 -250
rect 658 -286 666 -269
rect 1050 -286 1058 -269
rect 658 -294 1058 -286
rect 1087 -269 1487 -250
rect 1087 -286 1095 -269
rect 1479 -286 1487 -269
rect 1087 -294 1487 -286
<< polycont >>
rect -1479 269 -1095 286
rect -1050 269 -666 286
rect -621 269 -237 286
rect -192 269 192 286
rect 237 269 621 286
rect 666 269 1050 286
rect 1095 269 1479 286
rect -1479 -286 -1095 -269
rect -1050 -286 -666 -269
rect -621 -286 -237 -269
rect -192 -286 192 -269
rect 237 -286 621 -269
rect 666 -286 1050 -269
rect 1095 -286 1479 -269
<< locali >>
rect -1577 338 -1529 355
rect 1529 338 1577 355
rect -1577 307 -1560 338
rect 1560 307 1577 338
rect -1487 269 -1479 286
rect -1095 269 -1087 286
rect -1058 269 -1050 286
rect -666 269 -658 286
rect -629 269 -621 286
rect -237 269 -229 286
rect -200 269 -192 286
rect 192 269 200 286
rect 229 269 237 286
rect 621 269 629 286
rect 658 269 666 286
rect 1050 269 1058 286
rect 1087 269 1095 286
rect 1479 269 1487 286
rect -1510 244 -1493 252
rect -1510 -252 -1493 -244
rect -1081 244 -1064 252
rect -1081 -252 -1064 -244
rect -652 244 -635 252
rect -652 -252 -635 -244
rect -223 244 -206 252
rect -223 -252 -206 -244
rect 206 244 223 252
rect 206 -252 223 -244
rect 635 244 652 252
rect 635 -252 652 -244
rect 1064 244 1081 252
rect 1064 -252 1081 -244
rect 1493 244 1510 252
rect 1493 -252 1510 -244
rect -1487 -286 -1479 -269
rect -1095 -286 -1087 -269
rect -1058 -286 -1050 -269
rect -666 -286 -658 -269
rect -629 -286 -621 -269
rect -237 -286 -229 -269
rect -200 -286 -192 -269
rect 192 -286 200 -269
rect 229 -286 237 -269
rect 621 -286 629 -269
rect 658 -286 666 -269
rect 1050 -286 1058 -269
rect 1087 -286 1095 -269
rect 1479 -286 1487 -269
rect -1577 -338 -1560 -307
rect 1560 -338 1577 -307
rect -1577 -355 -1529 -338
rect 1529 -355 1577 -338
<< viali >>
rect -1479 269 -1095 286
rect -1050 269 -666 286
rect -621 269 -237 286
rect -192 269 192 286
rect 237 269 621 286
rect 666 269 1050 286
rect 1095 269 1479 286
rect -1510 -244 -1493 244
rect -1081 -244 -1064 244
rect -652 -244 -635 244
rect -223 -244 -206 244
rect 206 -244 223 244
rect 635 -244 652 244
rect 1064 -244 1081 244
rect 1493 -244 1510 244
rect -1479 -286 -1095 -269
rect -1050 -286 -666 -269
rect -621 -286 -237 -269
rect -192 -286 192 -269
rect 237 -286 621 -269
rect 666 -286 1050 -269
rect 1095 -286 1479 -269
<< metal1 >>
rect -1485 286 -1089 289
rect -1485 269 -1479 286
rect -1095 269 -1089 286
rect -1485 266 -1089 269
rect -1056 286 -660 289
rect -1056 269 -1050 286
rect -666 269 -660 286
rect -1056 266 -660 269
rect -627 286 -231 289
rect -627 269 -621 286
rect -237 269 -231 286
rect -627 266 -231 269
rect -198 286 198 289
rect -198 269 -192 286
rect 192 269 198 286
rect -198 266 198 269
rect 231 286 627 289
rect 231 269 237 286
rect 621 269 627 286
rect 231 266 627 269
rect 660 286 1056 289
rect 660 269 666 286
rect 1050 269 1056 286
rect 660 266 1056 269
rect 1089 286 1485 289
rect 1089 269 1095 286
rect 1479 269 1485 286
rect 1089 266 1485 269
rect -1513 244 -1490 250
rect -1513 -244 -1510 244
rect -1493 -244 -1490 244
rect -1513 -250 -1490 -244
rect -1084 244 -1061 250
rect -1084 -244 -1081 244
rect -1064 -244 -1061 244
rect -1084 -250 -1061 -244
rect -655 244 -632 250
rect -655 -244 -652 244
rect -635 -244 -632 244
rect -655 -250 -632 -244
rect -226 244 -203 250
rect -226 -244 -223 244
rect -206 -244 -203 244
rect -226 -250 -203 -244
rect 203 244 226 250
rect 203 -244 206 244
rect 223 -244 226 244
rect 203 -250 226 -244
rect 632 244 655 250
rect 632 -244 635 244
rect 652 -244 655 244
rect 632 -250 655 -244
rect 1061 244 1084 250
rect 1061 -244 1064 244
rect 1081 -244 1084 244
rect 1061 -250 1084 -244
rect 1490 244 1513 250
rect 1490 -244 1493 244
rect 1510 -244 1513 244
rect 1490 -250 1513 -244
rect -1485 -269 -1089 -266
rect -1485 -286 -1479 -269
rect -1095 -286 -1089 -269
rect -1485 -289 -1089 -286
rect -1056 -269 -660 -266
rect -1056 -286 -1050 -269
rect -666 -286 -660 -269
rect -1056 -289 -660 -286
rect -627 -269 -231 -266
rect -627 -286 -621 -269
rect -237 -286 -231 -269
rect -627 -289 -231 -286
rect -198 -269 198 -266
rect -198 -286 -192 -269
rect 192 -286 198 -269
rect -198 -289 198 -286
rect 231 -269 627 -266
rect 231 -286 237 -269
rect 621 -286 627 -269
rect 231 -289 627 -286
rect 660 -269 1056 -266
rect 660 -286 666 -269
rect 1050 -286 1056 -269
rect 660 -289 1056 -286
rect 1089 -269 1485 -266
rect 1089 -286 1095 -269
rect 1479 -286 1485 -269
rect 1089 -289 1485 -286
<< properties >>
string FIXED_BBOX -1568 -346 1568 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 4 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
