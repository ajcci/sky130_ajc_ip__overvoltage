magic
tech sky130A
magscale 1 2
timestamp 1712066688
<< pwell >>
rect -3631 -758 3631 758
<< mvnmos >>
rect -3403 -500 -2603 500
rect -2545 -500 -1745 500
rect -1687 -500 -887 500
rect -829 -500 -29 500
rect 29 -500 829 500
rect 887 -500 1687 500
rect 1745 -500 2545 500
rect 2603 -500 3403 500
<< mvndiff >>
rect -3461 488 -3403 500
rect -3461 -488 -3449 488
rect -3415 -488 -3403 488
rect -3461 -500 -3403 -488
rect -2603 488 -2545 500
rect -2603 -488 -2591 488
rect -2557 -488 -2545 488
rect -2603 -500 -2545 -488
rect -1745 488 -1687 500
rect -1745 -488 -1733 488
rect -1699 -488 -1687 488
rect -1745 -500 -1687 -488
rect -887 488 -829 500
rect -887 -488 -875 488
rect -841 -488 -829 488
rect -887 -500 -829 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 829 488 887 500
rect 829 -488 841 488
rect 875 -488 887 488
rect 829 -500 887 -488
rect 1687 488 1745 500
rect 1687 -488 1699 488
rect 1733 -488 1745 488
rect 1687 -500 1745 -488
rect 2545 488 2603 500
rect 2545 -488 2557 488
rect 2591 -488 2603 488
rect 2545 -500 2603 -488
rect 3403 488 3461 500
rect 3403 -488 3415 488
rect 3449 -488 3461 488
rect 3403 -500 3461 -488
<< mvndiffc >>
rect -3449 -488 -3415 488
rect -2591 -488 -2557 488
rect -1733 -488 -1699 488
rect -875 -488 -841 488
rect -17 -488 17 488
rect 841 -488 875 488
rect 1699 -488 1733 488
rect 2557 -488 2591 488
rect 3415 -488 3449 488
<< mvpsubdiff >>
rect -3595 710 3595 722
rect -3595 676 -3487 710
rect 3487 676 3595 710
rect -3595 664 3595 676
rect -3595 614 -3537 664
rect -3595 -614 -3583 614
rect -3549 -614 -3537 614
rect 3537 614 3595 664
rect -3595 -664 -3537 -614
rect 3537 -614 3549 614
rect 3583 -614 3595 614
rect 3537 -664 3595 -614
rect -3595 -676 3595 -664
rect -3595 -710 -3487 -676
rect 3487 -710 3595 -676
rect -3595 -722 3595 -710
<< mvpsubdiffcont >>
rect -3487 676 3487 710
rect -3583 -614 -3549 614
rect 3549 -614 3583 614
rect -3487 -710 3487 -676
<< poly >>
rect -3403 572 -2603 588
rect -3403 538 -3387 572
rect -2619 538 -2603 572
rect -3403 500 -2603 538
rect -2545 572 -1745 588
rect -2545 538 -2529 572
rect -1761 538 -1745 572
rect -2545 500 -1745 538
rect -1687 572 -887 588
rect -1687 538 -1671 572
rect -903 538 -887 572
rect -1687 500 -887 538
rect -829 572 -29 588
rect -829 538 -813 572
rect -45 538 -29 572
rect -829 500 -29 538
rect 29 572 829 588
rect 29 538 45 572
rect 813 538 829 572
rect 29 500 829 538
rect 887 572 1687 588
rect 887 538 903 572
rect 1671 538 1687 572
rect 887 500 1687 538
rect 1745 572 2545 588
rect 1745 538 1761 572
rect 2529 538 2545 572
rect 1745 500 2545 538
rect 2603 572 3403 588
rect 2603 538 2619 572
rect 3387 538 3403 572
rect 2603 500 3403 538
rect -3403 -538 -2603 -500
rect -3403 -572 -3387 -538
rect -2619 -572 -2603 -538
rect -3403 -588 -2603 -572
rect -2545 -538 -1745 -500
rect -2545 -572 -2529 -538
rect -1761 -572 -1745 -538
rect -2545 -588 -1745 -572
rect -1687 -538 -887 -500
rect -1687 -572 -1671 -538
rect -903 -572 -887 -538
rect -1687 -588 -887 -572
rect -829 -538 -29 -500
rect -829 -572 -813 -538
rect -45 -572 -29 -538
rect -829 -588 -29 -572
rect 29 -538 829 -500
rect 29 -572 45 -538
rect 813 -572 829 -538
rect 29 -588 829 -572
rect 887 -538 1687 -500
rect 887 -572 903 -538
rect 1671 -572 1687 -538
rect 887 -588 1687 -572
rect 1745 -538 2545 -500
rect 1745 -572 1761 -538
rect 2529 -572 2545 -538
rect 1745 -588 2545 -572
rect 2603 -538 3403 -500
rect 2603 -572 2619 -538
rect 3387 -572 3403 -538
rect 2603 -588 3403 -572
<< polycont >>
rect -3387 538 -2619 572
rect -2529 538 -1761 572
rect -1671 538 -903 572
rect -813 538 -45 572
rect 45 538 813 572
rect 903 538 1671 572
rect 1761 538 2529 572
rect 2619 538 3387 572
rect -3387 -572 -2619 -538
rect -2529 -572 -1761 -538
rect -1671 -572 -903 -538
rect -813 -572 -45 -538
rect 45 -572 813 -538
rect 903 -572 1671 -538
rect 1761 -572 2529 -538
rect 2619 -572 3387 -538
<< locali >>
rect -3583 676 -3487 710
rect 3487 676 3583 710
rect -3583 614 -3549 676
rect 3549 614 3583 676
rect -3403 538 -3387 572
rect -2619 538 -2603 572
rect -2545 538 -2529 572
rect -1761 538 -1745 572
rect -1687 538 -1671 572
rect -903 538 -887 572
rect -829 538 -813 572
rect -45 538 -29 572
rect 29 538 45 572
rect 813 538 829 572
rect 887 538 903 572
rect 1671 538 1687 572
rect 1745 538 1761 572
rect 2529 538 2545 572
rect 2603 538 2619 572
rect 3387 538 3403 572
rect -3449 488 -3415 504
rect -3449 -504 -3415 -488
rect -2591 488 -2557 504
rect -2591 -504 -2557 -488
rect -1733 488 -1699 504
rect -1733 -504 -1699 -488
rect -875 488 -841 504
rect -875 -504 -841 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 841 488 875 504
rect 841 -504 875 -488
rect 1699 488 1733 504
rect 1699 -504 1733 -488
rect 2557 488 2591 504
rect 2557 -504 2591 -488
rect 3415 488 3449 504
rect 3415 -504 3449 -488
rect -3403 -572 -3387 -538
rect -2619 -572 -2603 -538
rect -2545 -572 -2529 -538
rect -1761 -572 -1745 -538
rect -1687 -572 -1671 -538
rect -903 -572 -887 -538
rect -829 -572 -813 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 813 -572 829 -538
rect 887 -572 903 -538
rect 1671 -572 1687 -538
rect 1745 -572 1761 -538
rect 2529 -572 2545 -538
rect 2603 -572 2619 -538
rect 3387 -572 3403 -538
rect -3583 -676 -3549 -614
rect 3549 -676 3583 -614
rect -3583 -710 -3487 -676
rect 3487 -710 3583 -676
<< viali >>
rect -3387 538 -2619 572
rect -2529 538 -1761 572
rect -1671 538 -903 572
rect -813 538 -45 572
rect 45 538 813 572
rect 903 538 1671 572
rect 1761 538 2529 572
rect 2619 538 3387 572
rect -3449 -488 -3415 488
rect -2591 -488 -2557 488
rect -1733 -488 -1699 488
rect -875 -488 -841 488
rect -17 -488 17 488
rect 841 -488 875 488
rect 1699 -488 1733 488
rect 2557 -488 2591 488
rect 3415 -488 3449 488
rect -3387 -572 -2619 -538
rect -2529 -572 -1761 -538
rect -1671 -572 -903 -538
rect -813 -572 -45 -538
rect 45 -572 813 -538
rect 903 -572 1671 -538
rect 1761 -572 2529 -538
rect 2619 -572 3387 -538
<< metal1 >>
rect -3399 572 -2607 578
rect -3399 538 -3387 572
rect -2619 538 -2607 572
rect -3399 532 -2607 538
rect -2541 572 -1749 578
rect -2541 538 -2529 572
rect -1761 538 -1749 572
rect -2541 532 -1749 538
rect -1683 572 -891 578
rect -1683 538 -1671 572
rect -903 538 -891 572
rect -1683 532 -891 538
rect -825 572 -33 578
rect -825 538 -813 572
rect -45 538 -33 572
rect -825 532 -33 538
rect 33 572 825 578
rect 33 538 45 572
rect 813 538 825 572
rect 33 532 825 538
rect 891 572 1683 578
rect 891 538 903 572
rect 1671 538 1683 572
rect 891 532 1683 538
rect 1749 572 2541 578
rect 1749 538 1761 572
rect 2529 538 2541 572
rect 1749 532 2541 538
rect 2607 572 3399 578
rect 2607 538 2619 572
rect 3387 538 3399 572
rect 2607 532 3399 538
rect -3455 488 -3409 500
rect -3455 -488 -3449 488
rect -3415 -488 -3409 488
rect -3455 -500 -3409 -488
rect -2597 488 -2551 500
rect -2597 -488 -2591 488
rect -2557 -488 -2551 488
rect -2597 -500 -2551 -488
rect -1739 488 -1693 500
rect -1739 -488 -1733 488
rect -1699 -488 -1693 488
rect -1739 -500 -1693 -488
rect -881 488 -835 500
rect -881 -488 -875 488
rect -841 -488 -835 488
rect -881 -500 -835 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 835 488 881 500
rect 835 -488 841 488
rect 875 -488 881 488
rect 835 -500 881 -488
rect 1693 488 1739 500
rect 1693 -488 1699 488
rect 1733 -488 1739 488
rect 1693 -500 1739 -488
rect 2551 488 2597 500
rect 2551 -488 2557 488
rect 2591 -488 2597 488
rect 2551 -500 2597 -488
rect 3409 488 3455 500
rect 3409 -488 3415 488
rect 3449 -488 3455 488
rect 3409 -500 3455 -488
rect -3399 -538 -2607 -532
rect -3399 -572 -3387 -538
rect -2619 -572 -2607 -538
rect -3399 -578 -2607 -572
rect -2541 -538 -1749 -532
rect -2541 -572 -2529 -538
rect -1761 -572 -1749 -538
rect -2541 -578 -1749 -572
rect -1683 -538 -891 -532
rect -1683 -572 -1671 -538
rect -903 -572 -891 -538
rect -1683 -578 -891 -572
rect -825 -538 -33 -532
rect -825 -572 -813 -538
rect -45 -572 -33 -538
rect -825 -578 -33 -572
rect 33 -538 825 -532
rect 33 -572 45 -538
rect 813 -572 825 -538
rect 33 -578 825 -572
rect 891 -538 1683 -532
rect 891 -572 903 -538
rect 1671 -572 1683 -538
rect 891 -578 1683 -572
rect 1749 -538 2541 -532
rect 1749 -572 1761 -538
rect 2529 -572 2541 -538
rect 1749 -578 2541 -572
rect 2607 -538 3399 -532
rect 2607 -572 2619 -538
rect 3387 -572 3399 -538
rect 2607 -578 3399 -572
<< properties >>
string FIXED_BBOX -3566 -693 3566 693
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 4 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
