magic
tech sky130A
magscale 1 2
timestamp 1711636687
<< nwell >>
rect -1887 -347 1887 347
<< mvpmos >>
rect -1629 -50 -29 50
rect 29 -50 1629 50
<< mvpdiff >>
rect -1687 38 -1629 50
rect -1687 -38 -1675 38
rect -1641 -38 -1629 38
rect -1687 -50 -1629 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 1629 38 1687 50
rect 1629 -38 1641 38
rect 1675 -38 1687 38
rect 1629 -50 1687 -38
<< mvpdiffc >>
rect -1675 -38 -1641 38
rect -17 -38 17 38
rect 1641 -38 1675 38
<< mvnsubdiff >>
rect -1821 269 1821 281
rect -1821 235 -1713 269
rect 1713 235 1821 269
rect -1821 223 1821 235
rect -1821 173 -1763 223
rect -1821 -173 -1809 173
rect -1775 -173 -1763 173
rect 1763 173 1821 223
rect -1821 -223 -1763 -173
rect 1763 -173 1775 173
rect 1809 -173 1821 173
rect 1763 -223 1821 -173
rect -1821 -235 1821 -223
rect -1821 -269 -1713 -235
rect 1713 -269 1821 -235
rect -1821 -281 1821 -269
<< mvnsubdiffcont >>
rect -1713 235 1713 269
rect -1809 -173 -1775 173
rect 1775 -173 1809 173
rect -1713 -269 1713 -235
<< poly >>
rect -1629 131 -29 147
rect -1629 97 -1613 131
rect -45 97 -29 131
rect -1629 50 -29 97
rect 29 131 1629 147
rect 29 97 45 131
rect 1613 97 1629 131
rect 29 50 1629 97
rect -1629 -97 -29 -50
rect -1629 -131 -1613 -97
rect -45 -131 -29 -97
rect -1629 -147 -29 -131
rect 29 -97 1629 -50
rect 29 -131 45 -97
rect 1613 -131 1629 -97
rect 29 -147 1629 -131
<< polycont >>
rect -1613 97 -45 131
rect 45 97 1613 131
rect -1613 -131 -45 -97
rect 45 -131 1613 -97
<< locali >>
rect -1809 235 -1713 269
rect 1713 235 1809 269
rect -1809 173 -1775 235
rect 1775 173 1809 235
rect -1629 97 -1613 131
rect -45 97 -29 131
rect 29 97 45 131
rect 1613 97 1629 131
rect -1675 38 -1641 54
rect -1675 -54 -1641 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 1641 38 1675 54
rect 1641 -54 1675 -38
rect -1629 -131 -1613 -97
rect -45 -131 -29 -97
rect 29 -131 45 -97
rect 1613 -131 1629 -97
rect -1809 -235 -1775 -173
rect 1775 -235 1809 -173
rect -1809 -269 -1713 -235
rect 1713 -269 1809 -235
<< viali >>
rect -1613 97 -45 131
rect 45 97 1613 131
rect -1675 -38 -1641 38
rect -17 -38 17 38
rect 1641 -38 1675 38
rect -1613 -131 -45 -97
rect 45 -131 1613 -97
<< metal1 >>
rect -1625 131 -33 137
rect -1625 97 -1613 131
rect -45 97 -33 131
rect -1625 91 -33 97
rect 33 131 1625 137
rect 33 97 45 131
rect 1613 97 1625 131
rect 33 91 1625 97
rect -1681 38 -1635 50
rect -1681 -38 -1675 38
rect -1641 -38 -1635 38
rect -1681 -50 -1635 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 1635 38 1681 50
rect 1635 -38 1641 38
rect 1675 -38 1681 38
rect 1635 -50 1681 -38
rect -1625 -97 -33 -91
rect -1625 -131 -1613 -97
rect -45 -131 -33 -97
rect -1625 -137 -33 -131
rect 33 -97 1625 -91
rect 33 -131 45 -97
rect 1613 -131 1625 -97
rect 33 -137 1625 -131
<< properties >>
string FIXED_BBOX -1792 -252 1792 252
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 8.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
